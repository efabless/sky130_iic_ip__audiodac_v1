magic
tech sky130A
timestamp 1644659262
<< nwell >>
rect 917 -12717 1612 -11420
<< pwell >>
rect 932 -13501 1597 -12743
<< mvnmos >>
rect 1046 -13372 1096 -12872
rect 1125 -13372 1175 -12872
rect 1354 -13372 1404 -12872
rect 1433 -13372 1483 -12872
<< mvpmos >>
rect 1046 -12569 1096 -11569
rect 1125 -12569 1175 -11569
rect 1354 -12569 1404 -11569
rect 1433 -12569 1483 -11569
<< mvndiff >>
rect 1017 -12878 1046 -12872
rect 1017 -13366 1023 -12878
rect 1040 -13366 1046 -12878
rect 1017 -13372 1046 -13366
rect 1096 -12878 1125 -12872
rect 1096 -13366 1102 -12878
rect 1119 -13366 1125 -12878
rect 1096 -13372 1125 -13366
rect 1175 -12878 1204 -12872
rect 1175 -13366 1181 -12878
rect 1198 -13366 1204 -12878
rect 1175 -13372 1204 -13366
rect 1325 -12878 1354 -12872
rect 1325 -13366 1331 -12878
rect 1348 -13366 1354 -12878
rect 1325 -13372 1354 -13366
rect 1404 -12878 1433 -12872
rect 1404 -13366 1410 -12878
rect 1427 -13366 1433 -12878
rect 1404 -13372 1433 -13366
rect 1483 -12878 1512 -12872
rect 1483 -13366 1489 -12878
rect 1506 -13366 1512 -12878
rect 1483 -13372 1512 -13366
<< mvpdiff >>
rect 1017 -11575 1046 -11569
rect 1017 -12563 1023 -11575
rect 1040 -12563 1046 -11575
rect 1017 -12569 1046 -12563
rect 1096 -11575 1125 -11569
rect 1096 -12563 1102 -11575
rect 1119 -12563 1125 -11575
rect 1096 -12569 1125 -12563
rect 1175 -11575 1204 -11569
rect 1175 -12563 1181 -11575
rect 1198 -12563 1204 -11575
rect 1175 -12569 1204 -12563
rect 1325 -11575 1354 -11569
rect 1325 -12563 1331 -11575
rect 1348 -12563 1354 -11575
rect 1325 -12569 1354 -12563
rect 1404 -11575 1433 -11569
rect 1404 -12563 1410 -11575
rect 1427 -12563 1433 -11575
rect 1404 -12569 1433 -12563
rect 1483 -11575 1512 -11569
rect 1483 -12563 1489 -11575
rect 1506 -12563 1512 -11575
rect 1483 -12569 1512 -12563
<< mvndiffc >>
rect 1023 -13366 1040 -12878
rect 1102 -13366 1119 -12878
rect 1181 -13366 1198 -12878
rect 1331 -13366 1348 -12878
rect 1410 -13366 1427 -12878
rect 1489 -13366 1506 -12878
<< mvpdiffc >>
rect 1023 -12563 1040 -11575
rect 1102 -12563 1119 -11575
rect 1181 -12563 1198 -11575
rect 1331 -12563 1348 -11575
rect 1410 -12563 1427 -11575
rect 1489 -12563 1506 -11575
<< mvpsubdiff >>
rect 950 -12767 1579 -12761
rect 950 -12784 1004 -12767
rect 1217 -12784 1312 -12767
rect 1525 -12784 1579 -12767
rect 950 -12790 1579 -12784
rect 950 -12815 979 -12790
rect 950 -13429 956 -12815
rect 973 -13429 979 -12815
rect 1242 -12815 1287 -12790
rect 950 -13454 979 -13429
rect 1242 -13429 1248 -12815
rect 1281 -13429 1287 -12815
rect 1550 -12815 1579 -12790
rect 1242 -13454 1287 -13429
rect 1550 -13429 1556 -12815
rect 1573 -13429 1579 -12815
rect 1550 -13454 1579 -13429
rect 950 -13460 1579 -13454
rect 950 -13477 1004 -13460
rect 1217 -13477 1312 -13460
rect 1525 -13477 1579 -13460
rect 950 -13483 1579 -13477
<< mvnsubdiff >>
rect 950 -11459 1579 -11453
rect 950 -11476 1004 -11459
rect 1217 -11476 1312 -11459
rect 1525 -11476 1579 -11459
rect 950 -11482 1579 -11476
rect 950 -11507 979 -11482
rect 950 -12630 956 -11507
rect 973 -12630 979 -11507
rect 1242 -11507 1287 -11482
rect 950 -12655 979 -12630
rect 1242 -12630 1248 -11507
rect 1281 -12630 1287 -11507
rect 1550 -11507 1579 -11482
rect 1242 -12655 1287 -12630
rect 1550 -12630 1556 -11507
rect 1573 -12630 1579 -11507
rect 1550 -12655 1579 -12630
rect 950 -12661 1579 -12655
rect 950 -12678 1004 -12661
rect 1217 -12678 1312 -12661
rect 1525 -12678 1579 -12661
rect 950 -12684 1579 -12678
<< mvpsubdiffcont >>
rect 1004 -12784 1217 -12767
rect 1312 -12784 1525 -12767
rect 956 -13429 973 -12815
rect 1248 -13429 1281 -12815
rect 1556 -13429 1573 -12815
rect 1004 -13477 1217 -13460
rect 1312 -13477 1525 -13460
<< mvnsubdiffcont >>
rect 1004 -11476 1217 -11459
rect 1312 -11476 1525 -11459
rect 956 -12630 973 -11507
rect 1248 -12630 1281 -11507
rect 1556 -12630 1573 -11507
rect 1004 -12678 1217 -12661
rect 1312 -12678 1525 -12661
<< poly >>
rect 1046 -11528 1096 -11520
rect 1046 -11545 1054 -11528
rect 1088 -11545 1096 -11528
rect 1046 -11569 1096 -11545
rect 1125 -11528 1175 -11520
rect 1125 -11545 1133 -11528
rect 1167 -11545 1175 -11528
rect 1125 -11569 1175 -11545
rect 1046 -12593 1096 -12569
rect 1046 -12610 1054 -12593
rect 1088 -12610 1096 -12593
rect 1046 -12618 1096 -12610
rect 1125 -12593 1175 -12569
rect 1125 -12610 1133 -12593
rect 1167 -12610 1175 -12593
rect 1125 -12618 1175 -12610
rect 1354 -11528 1404 -11520
rect 1354 -11545 1362 -11528
rect 1396 -11545 1404 -11528
rect 1354 -11569 1404 -11545
rect 1433 -11528 1483 -11520
rect 1433 -11545 1441 -11528
rect 1475 -11545 1483 -11528
rect 1433 -11569 1483 -11545
rect 1354 -12593 1404 -12569
rect 1354 -12610 1362 -12593
rect 1396 -12610 1404 -12593
rect 1354 -12618 1404 -12610
rect 1433 -12593 1483 -12569
rect 1433 -12610 1441 -12593
rect 1475 -12610 1483 -12593
rect 1433 -12618 1483 -12610
rect 1046 -12836 1096 -12828
rect 1046 -12853 1054 -12836
rect 1088 -12853 1096 -12836
rect 1046 -12872 1096 -12853
rect 1125 -12836 1175 -12828
rect 1125 -12853 1133 -12836
rect 1167 -12853 1175 -12836
rect 1125 -12872 1175 -12853
rect 1046 -13391 1096 -13372
rect 1046 -13408 1054 -13391
rect 1088 -13408 1096 -13391
rect 1046 -13416 1096 -13408
rect 1125 -13391 1175 -13372
rect 1125 -13408 1133 -13391
rect 1167 -13408 1175 -13391
rect 1125 -13416 1175 -13408
rect 1354 -12836 1404 -12828
rect 1354 -12853 1362 -12836
rect 1396 -12853 1404 -12836
rect 1354 -12872 1404 -12853
rect 1433 -12836 1483 -12828
rect 1433 -12853 1441 -12836
rect 1475 -12853 1483 -12836
rect 1433 -12872 1483 -12853
rect 1354 -13391 1404 -13372
rect 1354 -13408 1362 -13391
rect 1396 -13408 1404 -13391
rect 1354 -13416 1404 -13408
rect 1433 -13391 1483 -13372
rect 1433 -13408 1441 -13391
rect 1475 -13408 1483 -13391
rect 1433 -13416 1483 -13408
<< polycont >>
rect 1054 -11545 1088 -11528
rect 1133 -11545 1167 -11528
rect 1054 -12610 1088 -12593
rect 1133 -12610 1167 -12593
rect 1362 -11545 1396 -11528
rect 1441 -11545 1475 -11528
rect 1362 -12610 1396 -12593
rect 1441 -12610 1475 -12593
rect 1054 -12853 1088 -12836
rect 1133 -12853 1167 -12836
rect 1054 -13408 1088 -13391
rect 1133 -13408 1167 -13391
rect 1362 -12853 1396 -12836
rect 1441 -12853 1475 -12836
rect 1362 -13408 1396 -13391
rect 1441 -13408 1475 -13391
<< locali >>
rect 956 -11476 1004 -11459
rect 1217 -11476 1312 -11459
rect 1525 -11476 1573 -11459
rect 956 -11507 973 -11476
rect 1248 -11507 1281 -11476
rect 1046 -11545 1054 -11528
rect 1088 -11545 1096 -11528
rect 1125 -11545 1133 -11528
rect 1167 -11545 1175 -11528
rect 1023 -11575 1040 -11567
rect 1023 -12571 1040 -12563
rect 1102 -11575 1119 -11567
rect 1102 -12571 1119 -12563
rect 1181 -11575 1198 -11567
rect 1556 -11507 1573 -11476
rect 1354 -11545 1362 -11528
rect 1396 -11545 1404 -11528
rect 1433 -11545 1441 -11528
rect 1475 -11545 1483 -11528
rect 1331 -11575 1348 -11567
rect 1181 -12571 1198 -12563
rect 1046 -12610 1054 -12593
rect 1088 -12610 1096 -12593
rect 1125 -12610 1133 -12593
rect 1167 -12610 1175 -12593
rect 956 -12661 973 -12630
rect 1331 -12571 1348 -12563
rect 1410 -11575 1427 -11567
rect 1410 -12571 1427 -12563
rect 1489 -11575 1506 -11567
rect 1489 -12571 1506 -12563
rect 1354 -12610 1362 -12593
rect 1396 -12610 1404 -12593
rect 1433 -12610 1441 -12593
rect 1475 -12610 1483 -12593
rect 1248 -12661 1281 -12630
rect 1556 -12661 1573 -12630
rect 956 -12678 1004 -12661
rect 1217 -12678 1312 -12661
rect 1525 -12678 1573 -12661
rect 956 -12784 1004 -12767
rect 1217 -12784 1312 -12767
rect 1525 -12784 1573 -12767
rect 956 -12815 973 -12784
rect 1248 -12815 1281 -12784
rect 1046 -12853 1054 -12836
rect 1088 -12853 1096 -12836
rect 1125 -12853 1133 -12836
rect 1167 -12853 1175 -12836
rect 1023 -12878 1040 -12870
rect 1023 -13374 1040 -13366
rect 1102 -12878 1119 -12870
rect 1102 -13374 1119 -13366
rect 1181 -12878 1198 -12870
rect 1556 -12815 1573 -12784
rect 1354 -12853 1362 -12836
rect 1396 -12853 1404 -12836
rect 1433 -12853 1441 -12836
rect 1475 -12853 1483 -12836
rect 1331 -12878 1348 -12870
rect 1181 -13374 1198 -13366
rect 1046 -13408 1054 -13391
rect 1088 -13408 1096 -13391
rect 1125 -13408 1133 -13391
rect 1167 -13408 1175 -13391
rect 956 -13460 973 -13429
rect 1331 -13374 1348 -13366
rect 1410 -12878 1427 -12870
rect 1410 -13374 1427 -13366
rect 1489 -12878 1506 -12870
rect 1489 -13374 1506 -13366
rect 1354 -13408 1362 -13391
rect 1396 -13408 1404 -13391
rect 1433 -13408 1441 -13391
rect 1475 -13408 1483 -13391
rect 1248 -13460 1281 -13429
rect 1556 -13460 1573 -13429
rect 956 -13477 1004 -13460
rect 1217 -13477 1312 -13460
rect 1525 -13477 1573 -13460
<< viali >>
rect 1054 -11545 1088 -11528
rect 1133 -11545 1167 -11528
rect 1023 -12563 1040 -11575
rect 1102 -12563 1119 -11575
rect 1181 -12563 1198 -11575
rect 1362 -11545 1396 -11528
rect 1441 -11545 1475 -11528
rect 1244 -11661 1248 -11576
rect 1248 -11661 1281 -11576
rect 1281 -11661 1286 -11576
rect 1054 -12610 1088 -12593
rect 1133 -12610 1167 -12593
rect 1331 -12563 1348 -11575
rect 1410 -12563 1427 -11575
rect 1489 -12563 1506 -11575
rect 1362 -12610 1396 -12593
rect 1441 -12610 1475 -12593
rect 1054 -12853 1088 -12836
rect 1133 -12853 1167 -12836
rect 1023 -13366 1040 -12878
rect 1102 -13366 1119 -12878
rect 1181 -13366 1198 -12878
rect 1362 -12853 1396 -12836
rect 1441 -12853 1475 -12836
rect 1243 -13353 1248 -13268
rect 1248 -13353 1281 -13268
rect 1281 -13353 1285 -13268
rect 1054 -13408 1088 -13391
rect 1133 -13408 1167 -13391
rect 1331 -13366 1348 -12878
rect 1410 -13366 1427 -12878
rect 1489 -13366 1506 -12878
rect 1362 -13408 1396 -13391
rect 1441 -13408 1475 -13391
<< metal1 >>
rect 1048 -11528 1094 -11525
rect 1048 -11545 1054 -11528
rect 1088 -11545 1094 -11528
rect 1048 -11548 1094 -11545
rect 1127 -11528 1173 -11525
rect 1127 -11545 1133 -11528
rect 1167 -11545 1173 -11528
rect 1127 -11548 1173 -11545
rect 1356 -11528 1402 -11525
rect 1356 -11545 1362 -11528
rect 1396 -11545 1402 -11528
rect 1356 -11548 1402 -11545
rect 1435 -11528 1481 -11525
rect 1435 -11545 1441 -11528
rect 1475 -11545 1481 -11528
rect 1435 -11548 1481 -11545
rect 1020 -11575 1043 -11569
rect 1020 -11576 1023 -11575
rect 1040 -11576 1043 -11575
rect 1099 -11575 1122 -11569
rect 1014 -11661 1019 -11576
rect 1045 -11661 1050 -11576
rect 1020 -12563 1023 -11661
rect 1040 -12563 1043 -11661
rect 1099 -12509 1102 -11575
rect 1119 -12509 1122 -11575
rect 1178 -11575 1201 -11569
rect 1178 -11576 1181 -11575
rect 1198 -11576 1201 -11575
rect 1241 -11576 1289 -11570
rect 1328 -11575 1351 -11569
rect 1328 -11576 1331 -11575
rect 1348 -11576 1351 -11575
rect 1407 -11575 1430 -11569
rect 1172 -11661 1177 -11576
rect 1203 -11661 1208 -11576
rect 1239 -11661 1244 -11576
rect 1286 -11661 1291 -11576
rect 1322 -11661 1327 -11576
rect 1353 -11661 1358 -11576
rect 1090 -12558 1095 -12509
rect 1128 -12558 1133 -12509
rect 1020 -12569 1043 -12563
rect 1099 -12563 1102 -12558
rect 1119 -12563 1122 -12558
rect 1099 -12569 1122 -12563
rect 1178 -12563 1181 -11661
rect 1198 -12563 1201 -11661
rect 1241 -11667 1289 -11661
rect 1178 -12569 1201 -12563
rect 1328 -12563 1331 -11661
rect 1348 -12563 1351 -11661
rect 1407 -12509 1410 -11575
rect 1427 -12509 1430 -11575
rect 1486 -11575 1509 -11569
rect 1486 -11576 1489 -11575
rect 1506 -11576 1509 -11575
rect 1480 -11661 1485 -11576
rect 1511 -11661 1516 -11576
rect 1397 -12558 1402 -12509
rect 1435 -12558 1440 -12509
rect 1328 -12569 1351 -12563
rect 1407 -12563 1410 -12558
rect 1427 -12563 1430 -12558
rect 1407 -12569 1430 -12563
rect 1486 -12563 1489 -11661
rect 1506 -12563 1509 -11661
rect 1486 -12569 1509 -12563
rect 1048 -12593 1174 -12590
rect 1048 -12610 1054 -12593
rect 1088 -12610 1133 -12593
rect 1167 -12610 1174 -12593
rect 1048 -12758 1174 -12610
rect 1356 -12593 1482 -12590
rect 1356 -12610 1362 -12593
rect 1396 -12610 1441 -12593
rect 1475 -12610 1482 -12593
rect 1240 -12651 1289 -12648
rect 1356 -12651 1482 -12610
rect 1289 -12684 1482 -12651
rect 1240 -12687 1289 -12684
rect 1240 -12758 1289 -12755
rect 1048 -12791 1240 -12758
rect 1048 -12836 1174 -12791
rect 1240 -12794 1289 -12791
rect 1048 -12853 1054 -12836
rect 1088 -12853 1133 -12836
rect 1167 -12853 1174 -12836
rect 1048 -12856 1174 -12853
rect 1356 -12836 1482 -12684
rect 1356 -12853 1362 -12836
rect 1396 -12853 1441 -12836
rect 1475 -12853 1482 -12836
rect 1356 -12856 1482 -12853
rect 1020 -12878 1043 -12872
rect 1020 -13268 1023 -12878
rect 1040 -13268 1043 -12878
rect 1090 -12919 1095 -12870
rect 1128 -12919 1133 -12870
rect 1178 -12878 1201 -12872
rect 1014 -13353 1019 -13268
rect 1045 -13353 1050 -13268
rect 1020 -13366 1023 -13353
rect 1040 -13366 1043 -13353
rect 1020 -13372 1043 -13366
rect 1099 -13366 1102 -12919
rect 1119 -13366 1122 -12919
rect 1178 -13268 1181 -12878
rect 1198 -13268 1201 -12878
rect 1328 -12878 1351 -12872
rect 1240 -13268 1288 -13262
rect 1328 -13268 1331 -12878
rect 1348 -13268 1351 -12878
rect 1397 -12919 1402 -12870
rect 1435 -12919 1440 -12870
rect 1486 -12878 1509 -12872
rect 1172 -13353 1177 -13268
rect 1203 -13353 1208 -13268
rect 1238 -13353 1243 -13268
rect 1285 -13353 1290 -13268
rect 1322 -13353 1327 -13268
rect 1353 -13353 1358 -13268
rect 1099 -13372 1122 -13366
rect 1178 -13366 1181 -13353
rect 1198 -13366 1201 -13353
rect 1240 -13359 1288 -13353
rect 1178 -13372 1201 -13366
rect 1328 -13366 1331 -13353
rect 1348 -13366 1351 -13353
rect 1328 -13372 1351 -13366
rect 1407 -13366 1410 -12919
rect 1427 -13366 1430 -12919
rect 1486 -13268 1489 -12878
rect 1506 -13268 1509 -12878
rect 1479 -13353 1484 -13268
rect 1510 -13353 1515 -13268
rect 1407 -13372 1430 -13366
rect 1486 -13366 1489 -13353
rect 1506 -13366 1509 -13353
rect 1486 -13372 1509 -13366
rect 1048 -13391 1094 -13388
rect 1048 -13408 1054 -13391
rect 1088 -13408 1094 -13391
rect 1048 -13411 1094 -13408
rect 1127 -13391 1173 -13388
rect 1127 -13408 1133 -13391
rect 1167 -13408 1173 -13391
rect 1127 -13411 1173 -13408
rect 1356 -13391 1402 -13388
rect 1356 -13408 1362 -13391
rect 1396 -13408 1402 -13391
rect 1356 -13411 1402 -13408
rect 1435 -13391 1481 -13388
rect 1435 -13408 1441 -13391
rect 1475 -13408 1481 -13391
rect 1435 -13411 1481 -13408
<< via1 >>
rect 1019 -11661 1023 -11576
rect 1023 -11661 1040 -11576
rect 1040 -11661 1045 -11576
rect 1177 -11661 1181 -11576
rect 1181 -11661 1198 -11576
rect 1198 -11661 1203 -11576
rect 1244 -11661 1286 -11576
rect 1327 -11661 1331 -11576
rect 1331 -11661 1348 -11576
rect 1348 -11661 1353 -11576
rect 1095 -12558 1102 -12509
rect 1102 -12558 1119 -12509
rect 1119 -12558 1128 -12509
rect 1485 -11661 1489 -11576
rect 1489 -11661 1506 -11576
rect 1506 -11661 1511 -11576
rect 1402 -12558 1410 -12509
rect 1410 -12558 1427 -12509
rect 1427 -12558 1435 -12509
rect 1240 -12684 1289 -12651
rect 1240 -12791 1289 -12758
rect 1095 -12878 1128 -12870
rect 1095 -12919 1102 -12878
rect 1102 -12919 1119 -12878
rect 1119 -12919 1128 -12878
rect 1019 -13353 1023 -13268
rect 1023 -13353 1040 -13268
rect 1040 -13353 1045 -13268
rect 1402 -12878 1435 -12870
rect 1402 -12919 1410 -12878
rect 1410 -12919 1427 -12878
rect 1427 -12919 1435 -12878
rect 1177 -13353 1181 -13268
rect 1181 -13353 1198 -13268
rect 1198 -13353 1203 -13268
rect 1243 -13353 1285 -13268
rect 1327 -13353 1331 -13268
rect 1331 -13353 1348 -13268
rect 1348 -13353 1353 -13268
rect 1484 -13353 1489 -13268
rect 1489 -13353 1506 -13268
rect 1506 -13353 1510 -13268
<< metal2 >>
rect 1019 -11576 1045 -11571
rect 1177 -11576 1203 -11571
rect 1244 -11576 1286 -11571
rect 1327 -11576 1353 -11571
rect 1485 -11576 1511 -11571
rect 1045 -11661 1177 -11576
rect 1203 -11661 1244 -11576
rect 1286 -11661 1327 -11576
rect 1353 -11661 1485 -11576
rect 1019 -11666 1045 -11661
rect 1177 -11666 1203 -11661
rect 1244 -11666 1286 -11661
rect 1327 -11666 1353 -11661
rect 1485 -11666 1511 -11661
rect 1095 -12509 1128 -12504
rect 1095 -12651 1128 -12558
rect 1402 -12509 1435 -12504
rect 1095 -12684 1240 -12651
rect 1289 -12684 1292 -12651
rect 1095 -12870 1128 -12684
rect 1402 -12758 1435 -12558
rect 1237 -12791 1240 -12758
rect 1289 -12791 1435 -12758
rect 1095 -12924 1128 -12919
rect 1402 -12870 1435 -12791
rect 1402 -12924 1435 -12919
rect 1019 -13268 1045 -13263
rect 1177 -13268 1203 -13263
rect 1243 -13268 1285 -13263
rect 1327 -13268 1353 -13263
rect 1484 -13268 1510 -13263
rect 1045 -13353 1177 -13268
rect 1203 -13353 1243 -13268
rect 1285 -13353 1327 -13268
rect 1353 -13353 1484 -13268
rect 1019 -13358 1045 -13353
rect 1177 -13358 1203 -13353
rect 1243 -13358 1285 -13353
rect 1327 -13358 1353 -13353
rect 1484 -13358 1510 -13353
<< labels >>
rlabel metal2 1402 -12870 1435 -12558 1 in_n
port 2 n
rlabel metal2 1095 -12870 1128 -12558 1 in_p
port 1 n
rlabel metal2 1045 -13353 1177 -13268 1 vss
port 4 n
rlabel metal2 1045 -11661 1177 -11576 1 vdd_hi
port 3 n
<< end >>
