magic
tech sky130A
magscale 1 2
timestamp 1644660203
<< nwell >>
rect -4406 -7280 -3438 -7276
rect -4688 -8508 -3082 -7280
rect -4688 -8588 -3054 -8508
rect -4532 -9608 -3054 -8588
rect -4558 -10622 -2972 -9608
rect -4364 -11930 -3372 -10622
rect -4490 -13308 -3188 -11930
rect -4330 -14618 -3338 -13308
rect -3864 -15086 -3386 -14618
<< locali >>
rect -3960 -7376 -3764 -7354
rect -1922 -7376 -1778 -7354
rect 54 -7376 198 -7354
rect 2012 -7376 2156 -7354
rect 3974 -7376 4118 -7354
rect -3960 -7448 5946 -7376
rect -3960 -12004 -3764 -7448
rect -5572 -12128 -3764 -12004
rect -4980 -13324 -4850 -12128
rect -5572 -13380 -4850 -13324
rect -5572 -13514 -4856 -13380
rect -4978 -14058 -4866 -13514
rect -3960 -14546 -3764 -12128
rect -1922 -11114 -1778 -7448
rect -1922 -11598 -1920 -11114
rect -1782 -11598 -1778 -11114
rect -4890 -14805 -4271 -14799
rect -4890 -14867 -4884 -14805
rect -4822 -14867 -4271 -14805
rect -4890 -14873 -4271 -14867
rect -5078 -15278 -4952 -15178
rect -5510 -15322 -4952 -15278
rect -5510 -15408 -4954 -15322
rect -5070 -16582 -4954 -15408
rect -1922 -15552 -1778 -11598
rect -1786 -16036 -1778 -15552
rect -1922 -16410 -1778 -16036
rect 54 -8886 198 -7448
rect 54 -9370 60 -8886
rect 54 -13364 198 -9370
rect 54 -13848 58 -13364
rect 196 -13848 198 -13364
rect 54 -16410 198 -13848
rect 2012 -11114 2156 -7448
rect 3974 -8878 4118 -7448
rect 4110 -9362 4118 -8878
rect 2012 -11598 2016 -11114
rect 2154 -11598 2156 -11114
rect 2012 -15560 2156 -11598
rect 3974 -13368 4118 -9362
rect 4112 -13852 4118 -13368
rect 2012 -16044 2022 -15560
rect 2012 -16410 2156 -16044
rect 3974 -16410 4118 -13852
rect -3772 -16482 5966 -16410
rect -1922 -16500 -1778 -16482
rect 54 -16500 198 -16482
rect 2012 -16500 2156 -16482
rect 3974 -16500 4118 -16482
rect -5510 -16700 -3760 -16582
rect -1920 -16700 -1778 -16676
rect 54 -16700 196 -16676
rect 2014 -16700 2156 -16676
rect 3974 -16700 4116 -16676
rect -5510 -16706 5978 -16700
rect -3956 -18900 -3768 -16706
rect -3760 -16772 5978 -16706
rect -3960 -19000 -3768 -18900
rect -3960 -19102 -3774 -19000
rect -1920 -20390 -1778 -16772
rect -1920 -20874 -1918 -20390
rect -1780 -20874 -1778 -20390
rect -1920 -21220 -1778 -20874
rect 54 -18164 196 -16772
rect 54 -18648 56 -18164
rect 194 -18648 196 -18164
rect 54 -21220 196 -18648
rect 2014 -20388 2156 -16772
rect 3974 -18164 4116 -16772
rect 4110 -18648 4116 -18164
rect 2014 -20872 2016 -20388
rect 2154 -20872 2156 -20388
rect 2014 -21220 2156 -20872
rect 3974 -21220 4116 -18648
rect -3768 -21292 5970 -21220
rect -1920 -21314 -1778 -21292
rect 54 -21314 196 -21292
rect 2014 -21314 2156 -21292
rect 3974 -21314 4116 -21292
<< viali >>
rect -1920 -11598 -1782 -11114
rect -4884 -14867 -4822 -14805
rect -4271 -14873 -4197 -14799
rect -1924 -16036 -1786 -15552
rect 60 -9370 198 -8886
rect 58 -13848 196 -13364
rect 3972 -9362 4110 -8878
rect 2016 -11598 2154 -11114
rect 3974 -13852 4112 -13368
rect 2022 -16044 2160 -15560
rect -1918 -20874 -1780 -20390
rect 56 -18648 194 -18164
rect 3972 -18648 4110 -18164
rect 2016 -20872 2154 -20388
<< metal1 >>
rect -5708 -7798 -5698 -7668
rect -5638 -7798 -5628 -7668
rect -5396 -7796 -5386 -7666
rect -5326 -7796 -5316 -7666
rect -5076 -7798 -5066 -7668
rect -5006 -7798 -4996 -7668
rect -4762 -7796 -4752 -7666
rect -4692 -7796 -4682 -7666
rect -4446 -7798 -4436 -7668
rect -4376 -7798 -4366 -7668
rect -4130 -7798 -4120 -7668
rect -4060 -7798 -4050 -7668
rect -3554 -8536 -3544 -7666
rect -3418 -8536 -3408 -7666
rect -3236 -8536 -3226 -7666
rect -3100 -8536 -3090 -7666
rect -2922 -8538 -2912 -7668
rect -2786 -8538 -2776 -7668
rect -2606 -8538 -2596 -7668
rect -2470 -8538 -2460 -7668
rect -2288 -8538 -2278 -7668
rect -2152 -8538 -2142 -7668
rect -1568 -8536 -1558 -7666
rect -1432 -8536 -1422 -7666
rect -1250 -8536 -1240 -7666
rect -1114 -8536 -1104 -7666
rect -936 -8538 -926 -7668
rect -800 -8538 -790 -7668
rect -620 -8538 -610 -7668
rect -484 -8538 -474 -7668
rect -302 -8538 -292 -7668
rect -166 -8538 -156 -7668
rect 394 -8536 404 -7666
rect 530 -8536 540 -7666
rect 712 -8536 722 -7666
rect 848 -8536 858 -7666
rect 1026 -8538 1036 -7668
rect 1162 -8538 1172 -7668
rect 1342 -8538 1352 -7668
rect 1478 -8538 1488 -7668
rect 1660 -8538 1670 -7668
rect 1796 -8538 1806 -7668
rect 2356 -8542 2366 -7672
rect 2492 -8542 2502 -7672
rect 2674 -8542 2684 -7672
rect 2810 -8542 2820 -7672
rect 2988 -8544 2998 -7674
rect 3124 -8544 3134 -7674
rect 3304 -8544 3314 -7674
rect 3440 -8544 3450 -7674
rect 3622 -8544 3632 -7674
rect 3758 -8544 3768 -7674
rect 4314 -8542 4324 -7672
rect 4450 -8542 4460 -7672
rect 4632 -8542 4642 -7672
rect 4768 -8542 4778 -7672
rect 4946 -8544 4956 -7674
rect 5082 -8544 5092 -7674
rect 5262 -8544 5272 -7674
rect 5398 -8544 5408 -7674
rect 5580 -8544 5590 -7674
rect 5716 -8544 5726 -7674
rect -5554 -9500 -5544 -9370
rect -5484 -9500 -5474 -9370
rect -5236 -9500 -5226 -9370
rect -5166 -9500 -5156 -9370
rect -4920 -9500 -4910 -9370
rect -4850 -9500 -4840 -9370
rect -4608 -9502 -4598 -9372
rect -4538 -9502 -4528 -9372
rect -4292 -9502 -4282 -9372
rect -4222 -9502 -4212 -9372
rect -3708 -9524 -3698 -8654
rect -3572 -9524 -3562 -8654
rect -3390 -9524 -3380 -8654
rect -3254 -9524 -3244 -8654
rect -3076 -9526 -3066 -8656
rect -2940 -9526 -2930 -8656
rect -2760 -9526 -2750 -8656
rect -2624 -9526 -2614 -8656
rect -2442 -9526 -2432 -8656
rect -2306 -9526 -2296 -8656
rect -2128 -9526 -2118 -8656
rect -1992 -9526 -1982 -8656
rect -1722 -9524 -1712 -8654
rect -1586 -9524 -1576 -8654
rect -1404 -9524 -1394 -8654
rect -1268 -9524 -1258 -8654
rect -1090 -9526 -1080 -8656
rect -954 -9526 -944 -8656
rect -774 -9526 -764 -8656
rect -638 -9526 -628 -8656
rect -456 -9526 -446 -8656
rect -320 -9526 -310 -8656
rect -142 -9526 -132 -8656
rect -6 -9526 4 -8656
rect 54 -8886 204 -8874
rect 50 -9370 60 -8886
rect 198 -9370 208 -8886
rect 54 -9382 204 -9370
rect 240 -9524 250 -8654
rect 376 -9524 386 -8654
rect 558 -9524 568 -8654
rect 694 -9524 704 -8654
rect 872 -9526 882 -8656
rect 1008 -9526 1018 -8656
rect 1188 -9526 1198 -8656
rect 1324 -9526 1334 -8656
rect 1506 -9526 1516 -8656
rect 1642 -9526 1652 -8656
rect 1820 -9526 1830 -8656
rect 1956 -9526 1966 -8656
rect 2202 -9530 2212 -8660
rect 2338 -9530 2348 -8660
rect 2520 -9530 2530 -8660
rect 2656 -9530 2666 -8660
rect 2834 -9532 2844 -8662
rect 2970 -9532 2980 -8662
rect 3150 -9532 3160 -8662
rect 3286 -9532 3296 -8662
rect 3468 -9532 3478 -8662
rect 3604 -9532 3614 -8662
rect 3782 -9532 3792 -8662
rect 3918 -9532 3928 -8662
rect 3966 -8878 4116 -8866
rect 3962 -9362 3972 -8878
rect 4110 -9362 4120 -8878
rect 3966 -9374 4116 -9362
rect 4160 -9530 4170 -8660
rect 4296 -9530 4306 -8660
rect 4478 -9530 4488 -8660
rect 4614 -9530 4624 -8660
rect 4792 -9532 4802 -8662
rect 4928 -9532 4938 -8662
rect 5108 -9532 5118 -8662
rect 5244 -9532 5254 -8662
rect 5426 -9532 5436 -8662
rect 5562 -9532 5572 -8662
rect 5740 -9532 5750 -8662
rect 5876 -9532 5886 -8662
rect -5902 -9770 -4118 -9610
rect -3455 -9617 5782 -9616
rect -3923 -9626 5782 -9617
rect -5902 -14916 -5742 -9770
rect -5552 -10038 -5542 -9908
rect -5482 -10038 -5472 -9908
rect -5236 -10036 -5226 -9906
rect -5166 -10036 -5156 -9906
rect -4922 -10036 -4912 -9906
rect -4852 -10036 -4842 -9906
rect -4606 -10034 -4596 -9904
rect -4536 -10034 -4526 -9904
rect -4292 -10034 -4282 -9904
rect -4222 -10034 -4212 -9904
rect -3926 -9948 -3916 -9626
rect -3776 -9770 5782 -9626
rect -3776 -9771 -3455 -9770
rect -3776 -9948 -3766 -9771
rect -5712 -11678 -5702 -11548
rect -5642 -11678 -5632 -11548
rect -5396 -11676 -5386 -11546
rect -5326 -11676 -5316 -11546
rect -5082 -11678 -5072 -11548
rect -5012 -11678 -5002 -11548
rect -4762 -11680 -4752 -11550
rect -4692 -11680 -4682 -11550
rect -4446 -11680 -4436 -11550
rect -4376 -11680 -4366 -11550
rect -4130 -11680 -4120 -11550
rect -4060 -11680 -4050 -11550
rect -5458 -12580 -5448 -12450
rect -5388 -12580 -5378 -12450
rect -5146 -12580 -5136 -12450
rect -5076 -12580 -5066 -12450
rect -4764 -12572 -4754 -12442
rect -4694 -12572 -4684 -12442
rect -4446 -12578 -4436 -12448
rect -4376 -12578 -4366 -12448
rect -4134 -12578 -4124 -12448
rect -4064 -12578 -4054 -12448
rect -5302 -13056 -5292 -12926
rect -5232 -13056 -5222 -12926
rect -5906 -15120 -5896 -14916
rect -5756 -15120 -5742 -14916
rect -5902 -16668 -5742 -15120
rect -5612 -13218 -5122 -13166
rect -5612 -13536 -5560 -13218
rect -5612 -13588 -5082 -13536
rect -5612 -14964 -5560 -13588
rect -5450 -13670 -5398 -13588
rect -5464 -13800 -5454 -13670
rect -5394 -13800 -5384 -13670
rect -5302 -13798 -5292 -13668
rect -5232 -13798 -5222 -13668
rect -5134 -13672 -5082 -13588
rect -5146 -13802 -5136 -13672
rect -5076 -13802 -5066 -13672
rect -5328 -14860 -5220 -13880
rect -3923 -14088 -3769 -9948
rect -3554 -10772 -3544 -9902
rect -3418 -10772 -3408 -9902
rect -3236 -10772 -3226 -9902
rect -3100 -10772 -3090 -9902
rect -2922 -10774 -2912 -9904
rect -2786 -10774 -2776 -9904
rect -2606 -10774 -2596 -9904
rect -2470 -10774 -2460 -9904
rect -2288 -10774 -2278 -9904
rect -2152 -10774 -2142 -9904
rect -1568 -10772 -1558 -9902
rect -1432 -10772 -1422 -9902
rect -1250 -10772 -1240 -9902
rect -1114 -10772 -1104 -9902
rect -936 -10774 -926 -9904
rect -800 -10774 -790 -9904
rect -620 -10774 -610 -9904
rect -484 -10774 -474 -9904
rect -302 -10774 -292 -9904
rect -166 -10774 -156 -9904
rect 394 -10772 404 -9902
rect 530 -10772 540 -9902
rect 712 -10772 722 -9902
rect 848 -10772 858 -9902
rect 1026 -10774 1036 -9904
rect 1162 -10774 1172 -9904
rect 1342 -10774 1352 -9904
rect 1478 -10774 1488 -9904
rect 1660 -10774 1670 -9904
rect 1796 -10774 1806 -9904
rect 2356 -10778 2366 -9908
rect 2492 -10778 2502 -9908
rect 2674 -10778 2684 -9908
rect 2810 -10778 2820 -9908
rect 2988 -10780 2998 -9910
rect 3124 -10780 3134 -9910
rect 3304 -10780 3314 -9910
rect 3440 -10780 3450 -9910
rect 3622 -10780 3632 -9910
rect 3758 -10780 3768 -9910
rect 4314 -10778 4324 -9908
rect 4450 -10778 4460 -9908
rect 4632 -10778 4642 -9908
rect 4768 -10778 4778 -9908
rect 4946 -10780 4956 -9910
rect 5082 -10780 5092 -9910
rect 5262 -10780 5272 -9910
rect 5398 -10780 5408 -9910
rect 5580 -10780 5590 -9910
rect 5716 -10780 5726 -9910
rect -3708 -11760 -3698 -10890
rect -3572 -11760 -3562 -10890
rect -3390 -11760 -3380 -10890
rect -3254 -11760 -3244 -10890
rect -3076 -11762 -3066 -10892
rect -2940 -11762 -2930 -10892
rect -2760 -11762 -2750 -10892
rect -2624 -11762 -2614 -10892
rect -2442 -11762 -2432 -10892
rect -2306 -11762 -2296 -10892
rect -2128 -11762 -2118 -10892
rect -1992 -11762 -1982 -10892
rect -1926 -11114 -1776 -11102
rect -1930 -11598 -1920 -11114
rect -1782 -11598 -1772 -11114
rect -1926 -11610 -1776 -11598
rect -1722 -11760 -1712 -10890
rect -1586 -11760 -1576 -10890
rect -1404 -11760 -1394 -10890
rect -1268 -11760 -1258 -10890
rect -1090 -11762 -1080 -10892
rect -954 -11762 -944 -10892
rect -774 -11762 -764 -10892
rect -638 -11762 -628 -10892
rect -456 -11762 -446 -10892
rect -320 -11762 -310 -10892
rect -142 -11762 -132 -10892
rect -6 -11762 4 -10892
rect 240 -11760 250 -10890
rect 376 -11760 386 -10890
rect 558 -11760 568 -10890
rect 694 -11760 704 -10890
rect 872 -11762 882 -10892
rect 1008 -11762 1018 -10892
rect 1188 -11762 1198 -10892
rect 1324 -11762 1334 -10892
rect 1506 -11762 1516 -10892
rect 1642 -11762 1652 -10892
rect 1820 -11762 1830 -10892
rect 1956 -11762 1966 -10892
rect 2010 -11114 2160 -11102
rect 2006 -11598 2016 -11114
rect 2154 -11598 2164 -11114
rect 2010 -11610 2160 -11598
rect 2202 -11766 2212 -10896
rect 2338 -11766 2348 -10896
rect 2520 -11766 2530 -10896
rect 2656 -11766 2666 -10896
rect 2834 -11768 2844 -10898
rect 2970 -11768 2980 -10898
rect 3150 -11768 3160 -10898
rect 3286 -11768 3296 -10898
rect 3468 -11768 3478 -10898
rect 3604 -11768 3614 -10898
rect 3782 -11768 3792 -10898
rect 3918 -11768 3928 -10898
rect 4160 -11766 4170 -10896
rect 4296 -11766 4306 -10896
rect 4478 -11766 4488 -10896
rect 4614 -11766 4624 -10896
rect 4792 -11768 4802 -10898
rect 4928 -11768 4938 -10898
rect 5108 -11768 5118 -10898
rect 5244 -11768 5254 -10898
rect 5426 -11768 5436 -10898
rect 5562 -11768 5572 -10898
rect 5740 -11768 5750 -10898
rect 5876 -11768 5886 -10898
rect -3554 -13008 -3544 -12138
rect -3418 -13008 -3408 -12138
rect -3236 -13008 -3226 -12138
rect -3100 -13008 -3090 -12138
rect -2922 -13010 -2912 -12140
rect -2786 -13010 -2776 -12140
rect -2606 -13010 -2596 -12140
rect -2470 -13010 -2460 -12140
rect -2288 -13010 -2278 -12140
rect -2152 -13010 -2142 -12140
rect -1568 -13008 -1558 -12138
rect -1432 -13008 -1422 -12138
rect -1250 -13008 -1240 -12138
rect -1114 -13008 -1104 -12138
rect -936 -13010 -926 -12140
rect -800 -13010 -790 -12140
rect -620 -13010 -610 -12140
rect -484 -13010 -474 -12140
rect -302 -13010 -292 -12140
rect -166 -13010 -156 -12140
rect 394 -13008 404 -12138
rect 530 -13008 540 -12138
rect 712 -13008 722 -12138
rect 848 -13008 858 -12138
rect 1026 -13010 1036 -12140
rect 1162 -13010 1172 -12140
rect 1342 -13010 1352 -12140
rect 1478 -13010 1488 -12140
rect 1660 -13010 1670 -12140
rect 1796 -13010 1806 -12140
rect 2356 -13014 2366 -12144
rect 2492 -13014 2502 -12144
rect 2674 -13014 2684 -12144
rect 2810 -13014 2820 -12144
rect 2988 -13016 2998 -12146
rect 3124 -13016 3134 -12146
rect 3304 -13016 3314 -12146
rect 3440 -13016 3450 -12146
rect 3622 -13016 3632 -12146
rect 3758 -13016 3768 -12146
rect 4314 -13014 4324 -12144
rect 4450 -13014 4460 -12144
rect 4632 -13014 4642 -12144
rect 4768 -13014 4778 -12144
rect 4946 -13016 4956 -12146
rect 5082 -13016 5092 -12146
rect 5262 -13016 5272 -12146
rect 5398 -13016 5408 -12146
rect 5580 -13016 5590 -12146
rect 5716 -13016 5726 -12146
rect -3708 -13996 -3698 -13126
rect -3572 -13996 -3562 -13126
rect -3390 -13996 -3380 -13126
rect -3254 -13996 -3244 -13126
rect -3076 -13998 -3066 -13128
rect -2940 -13998 -2930 -13128
rect -2760 -13998 -2750 -13128
rect -2624 -13998 -2614 -13128
rect -2442 -13998 -2432 -13128
rect -2306 -13998 -2296 -13128
rect -2128 -13998 -2118 -13128
rect -1992 -13998 -1982 -13128
rect -1722 -13996 -1712 -13126
rect -1586 -13996 -1576 -13126
rect -1404 -13996 -1394 -13126
rect -1268 -13996 -1258 -13126
rect -1090 -13998 -1080 -13128
rect -954 -13998 -944 -13128
rect -774 -13998 -764 -13128
rect -638 -13998 -628 -13128
rect -456 -13998 -446 -13128
rect -320 -13998 -310 -13128
rect -142 -13998 -132 -13128
rect -6 -13998 4 -13128
rect 52 -13364 202 -13352
rect 48 -13848 58 -13364
rect 196 -13848 206 -13364
rect 52 -13860 202 -13848
rect 240 -13996 250 -13126
rect 376 -13996 386 -13126
rect 558 -13996 568 -13126
rect 694 -13996 704 -13126
rect 872 -13998 882 -13128
rect 1008 -13998 1018 -13128
rect 1188 -13998 1198 -13128
rect 1324 -13998 1334 -13128
rect 1506 -13998 1516 -13128
rect 1642 -13998 1652 -13128
rect 1820 -13998 1830 -13128
rect 1956 -13998 1966 -13128
rect 2202 -14002 2212 -13132
rect 2338 -14002 2348 -13132
rect 2520 -14002 2530 -13132
rect 2656 -14002 2666 -13132
rect 2834 -14004 2844 -13134
rect 2970 -14004 2980 -13134
rect 3150 -14004 3160 -13134
rect 3286 -14004 3296 -13134
rect 3468 -14004 3478 -13134
rect 3604 -14004 3614 -13134
rect 3782 -14004 3792 -13134
rect 3918 -14004 3928 -13134
rect 3968 -13368 4118 -13356
rect 3964 -13852 3974 -13368
rect 4112 -13852 4122 -13368
rect 3968 -13864 4118 -13852
rect 4160 -14002 4170 -13132
rect 4296 -14002 4306 -13132
rect 4478 -14002 4488 -13132
rect 4614 -14002 4624 -13132
rect 4792 -14004 4802 -13134
rect 4928 -14004 4938 -13134
rect 5108 -14004 5118 -13134
rect 5244 -14004 5254 -13134
rect 5426 -14004 5436 -13134
rect 5562 -14004 5572 -13134
rect 5740 -14004 5750 -13134
rect 5876 -14004 5886 -13134
rect -4604 -14248 -4594 -14118
rect -4534 -14248 -4524 -14118
rect -4284 -14246 -4274 -14116
rect -4214 -14246 -4204 -14116
rect -3923 -14242 5782 -14088
rect -4692 -14418 -4118 -14362
rect -4616 -14540 -4526 -14418
rect -4656 -14662 -4646 -14540
rect -4538 -14662 -4526 -14540
rect -4934 -14805 -4802 -14788
rect -4934 -14867 -4884 -14805
rect -4822 -14867 -4802 -14805
rect -4934 -14894 -4802 -14867
rect -5612 -15016 -5348 -14964
rect -5216 -14968 -4802 -14894
rect -5612 -15506 -5560 -15016
rect -4616 -15135 -4526 -14662
rect -4310 -14799 -4154 -14764
rect -4310 -14873 -4271 -14799
rect -4197 -14873 -4154 -14799
rect -4310 -14933 -4154 -14873
rect -4310 -15007 -4271 -14933
rect -4197 -15007 -4154 -14933
rect -4310 -15036 -4154 -15007
rect -5059 -15225 -4526 -15135
rect -5612 -15558 -5236 -15506
rect -5059 -15853 -4969 -15225
rect -4616 -15304 -4526 -15225
rect -4794 -15360 -4220 -15304
rect -4704 -15624 -4694 -15494
rect -4634 -15624 -4624 -15494
rect -4386 -15624 -4376 -15494
rect -4316 -15624 -4306 -15494
rect -5205 -15943 -4969 -15853
rect -5410 -16318 -5400 -16184
rect -5330 -16318 -5320 -16184
rect -4860 -16316 -4850 -16186
rect -4790 -16316 -4780 -16186
rect -4540 -16314 -4530 -16184
rect -4470 -16314 -4460 -16184
rect -4230 -16320 -4220 -16190
rect -4160 -16320 -4150 -16190
rect -5902 -16802 -4124 -16668
rect -5902 -16858 -4122 -16802
rect -3923 -16912 -3769 -14242
rect -3554 -15244 -3544 -14374
rect -3418 -15244 -3408 -14374
rect -3236 -15244 -3226 -14374
rect -3100 -15244 -3090 -14374
rect -2922 -15246 -2912 -14376
rect -2786 -15246 -2776 -14376
rect -2606 -15246 -2596 -14376
rect -2470 -15246 -2460 -14376
rect -2288 -15246 -2278 -14376
rect -2152 -15246 -2142 -14376
rect -1568 -15244 -1558 -14374
rect -1432 -15244 -1422 -14374
rect -1250 -15244 -1240 -14374
rect -1114 -15244 -1104 -14374
rect -936 -15246 -926 -14376
rect -800 -15246 -790 -14376
rect -620 -15246 -610 -14376
rect -484 -15246 -474 -14376
rect -302 -15246 -292 -14376
rect -166 -15246 -156 -14376
rect 394 -15244 404 -14374
rect 530 -15244 540 -14374
rect 712 -15244 722 -14374
rect 848 -15244 858 -14374
rect 1026 -15246 1036 -14376
rect 1162 -15246 1172 -14376
rect 1342 -15246 1352 -14376
rect 1478 -15246 1488 -14376
rect 1660 -15246 1670 -14376
rect 1796 -15246 1806 -14376
rect 2356 -15250 2366 -14380
rect 2492 -15250 2502 -14380
rect 2674 -15250 2684 -14380
rect 2810 -15250 2820 -14380
rect 2988 -15252 2998 -14382
rect 3124 -15252 3134 -14382
rect 3304 -15252 3314 -14382
rect 3440 -15252 3450 -14382
rect 3622 -15252 3632 -14382
rect 3758 -15252 3768 -14382
rect 4314 -15250 4324 -14380
rect 4450 -15250 4460 -14380
rect 4632 -15250 4642 -14380
rect 4768 -15250 4778 -14380
rect 4946 -15252 4956 -14382
rect 5082 -15252 5092 -14382
rect 5262 -15252 5272 -14382
rect 5398 -15252 5408 -14382
rect 5580 -15252 5590 -14382
rect 5716 -15252 5726 -14382
rect -3708 -16232 -3698 -15362
rect -3572 -16232 -3562 -15362
rect -3390 -16232 -3380 -15362
rect -3254 -16232 -3244 -15362
rect -3076 -16234 -3066 -15364
rect -2940 -16234 -2930 -15364
rect -2760 -16234 -2750 -15364
rect -2624 -16234 -2614 -15364
rect -2442 -16234 -2432 -15364
rect -2306 -16234 -2296 -15364
rect -2128 -16234 -2118 -15364
rect -1992 -16234 -1982 -15364
rect -1930 -15552 -1780 -15540
rect -1934 -16036 -1924 -15552
rect -1786 -16036 -1776 -15552
rect -1930 -16048 -1780 -16036
rect -1722 -16232 -1712 -15362
rect -1586 -16232 -1576 -15362
rect -1404 -16232 -1394 -15362
rect -1268 -16232 -1258 -15362
rect -1090 -16234 -1080 -15364
rect -954 -16234 -944 -15364
rect -774 -16234 -764 -15364
rect -638 -16234 -628 -15364
rect -456 -16234 -446 -15364
rect -320 -16234 -310 -15364
rect -142 -16234 -132 -15364
rect -6 -16234 4 -15364
rect 240 -16232 250 -15362
rect 376 -16232 386 -15362
rect 558 -16232 568 -15362
rect 694 -16232 704 -15362
rect 872 -16234 882 -15364
rect 1008 -16234 1018 -15364
rect 1188 -16234 1198 -15364
rect 1324 -16234 1334 -15364
rect 1506 -16234 1516 -15364
rect 1642 -16234 1652 -15364
rect 1820 -16234 1830 -15364
rect 1956 -16234 1966 -15364
rect 2016 -15560 2166 -15548
rect 2012 -16044 2022 -15560
rect 2160 -16044 2170 -15560
rect 2016 -16056 2166 -16044
rect 2202 -16238 2212 -15368
rect 2338 -16238 2348 -15368
rect 2520 -16238 2530 -15368
rect 2656 -16238 2666 -15368
rect 2834 -16240 2844 -15370
rect 2970 -16240 2980 -15370
rect 3150 -16240 3160 -15370
rect 3286 -16240 3296 -15370
rect 3468 -16240 3478 -15370
rect 3604 -16240 3614 -15370
rect 3782 -16240 3792 -15370
rect 3918 -16240 3928 -15370
rect 4160 -16238 4170 -15368
rect 4296 -16238 4306 -15368
rect 4478 -16238 4488 -15368
rect 4614 -16238 4624 -15368
rect 4792 -16240 4802 -15370
rect 4928 -16240 4938 -15370
rect 5108 -16240 5118 -15370
rect 5244 -16240 5254 -15370
rect 5426 -16240 5436 -15370
rect 5562 -16240 5572 -15370
rect 5740 -16240 5750 -15370
rect 5876 -16240 5886 -15370
rect -5552 -17124 -5542 -16994
rect -5482 -17124 -5472 -16994
rect -5238 -17124 -5228 -16994
rect -5168 -17124 -5158 -16994
rect -4922 -17126 -4912 -16996
rect -4852 -17126 -4842 -16996
rect -4604 -17126 -4594 -16996
rect -4534 -17126 -4524 -16996
rect -4286 -17128 -4276 -16998
rect -4216 -17128 -4206 -16998
rect -3923 -17170 -3908 -16912
rect -3786 -17170 -3769 -16912
rect -5712 -18774 -5702 -18644
rect -5642 -18774 -5632 -18644
rect -5396 -18776 -5386 -18646
rect -5326 -18776 -5316 -18646
rect -5078 -18776 -5068 -18646
rect -5008 -18776 -4998 -18646
rect -4762 -18776 -4752 -18646
rect -4692 -18776 -4682 -18646
rect -4446 -18776 -4436 -18646
rect -4376 -18776 -4366 -18646
rect -4128 -18776 -4118 -18646
rect -4058 -18776 -4048 -18646
rect -3923 -18920 -3769 -17170
rect -3554 -17850 -3544 -16980
rect -3418 -17850 -3408 -16980
rect -3236 -17850 -3226 -16980
rect -3100 -17850 -3090 -16980
rect -2922 -17852 -2912 -16982
rect -2786 -17852 -2776 -16982
rect -2606 -17852 -2596 -16982
rect -2470 -17852 -2460 -16982
rect -2288 -17852 -2278 -16982
rect -2152 -17852 -2142 -16982
rect -1568 -17850 -1558 -16980
rect -1432 -17850 -1422 -16980
rect -1250 -17850 -1240 -16980
rect -1114 -17850 -1104 -16980
rect -936 -17852 -926 -16982
rect -800 -17852 -790 -16982
rect -620 -17852 -610 -16982
rect -484 -17852 -474 -16982
rect -302 -17852 -292 -16982
rect -166 -17852 -156 -16982
rect 394 -17850 404 -16980
rect 530 -17850 540 -16980
rect 712 -17850 722 -16980
rect 848 -17850 858 -16980
rect 1026 -17852 1036 -16982
rect 1162 -17852 1172 -16982
rect 1342 -17852 1352 -16982
rect 1478 -17852 1488 -16982
rect 1660 -17852 1670 -16982
rect 1796 -17852 1806 -16982
rect 2356 -17856 2366 -16986
rect 2492 -17856 2502 -16986
rect 2674 -17856 2684 -16986
rect 2810 -17856 2820 -16986
rect 2988 -17858 2998 -16988
rect 3124 -17858 3134 -16988
rect 3304 -17858 3314 -16988
rect 3440 -17858 3450 -16988
rect 3622 -17858 3632 -16988
rect 3758 -17858 3768 -16988
rect 4314 -17856 4324 -16986
rect 4450 -17856 4460 -16986
rect 4632 -17856 4642 -16986
rect 4768 -17856 4778 -16986
rect 4946 -17858 4956 -16988
rect 5082 -17858 5092 -16988
rect 5262 -17858 5272 -16988
rect 5398 -17858 5408 -16988
rect 5580 -17858 5590 -16988
rect 5716 -17858 5726 -16988
rect -3708 -18838 -3698 -17968
rect -3572 -18838 -3562 -17968
rect -3390 -18838 -3380 -17968
rect -3254 -18838 -3244 -17968
rect -3076 -18840 -3066 -17970
rect -2940 -18840 -2930 -17970
rect -2760 -18840 -2750 -17970
rect -2624 -18840 -2614 -17970
rect -2442 -18840 -2432 -17970
rect -2306 -18840 -2296 -17970
rect -2128 -18840 -2118 -17970
rect -1992 -18840 -1982 -17970
rect -1722 -18838 -1712 -17968
rect -1586 -18838 -1576 -17968
rect -1404 -18838 -1394 -17968
rect -1268 -18838 -1258 -17968
rect -1090 -18840 -1080 -17970
rect -954 -18840 -944 -17970
rect -774 -18840 -764 -17970
rect -638 -18840 -628 -17970
rect -456 -18840 -446 -17970
rect -320 -18840 -310 -17970
rect -142 -18840 -132 -17970
rect -6 -18840 4 -17970
rect 50 -18164 200 -18152
rect 46 -18648 56 -18164
rect 194 -18648 204 -18164
rect 50 -18660 200 -18648
rect 240 -18838 250 -17968
rect 376 -18838 386 -17968
rect 558 -18838 568 -17968
rect 694 -18838 704 -17968
rect 872 -18840 882 -17970
rect 1008 -18840 1018 -17970
rect 1188 -18840 1198 -17970
rect 1324 -18840 1334 -17970
rect 1506 -18840 1516 -17970
rect 1642 -18840 1652 -17970
rect 1820 -18840 1830 -17970
rect 1956 -18840 1966 -17970
rect 2202 -18844 2212 -17974
rect 2338 -18844 2348 -17974
rect 2520 -18844 2530 -17974
rect 2656 -18844 2666 -17974
rect 2834 -18846 2844 -17976
rect 2970 -18846 2980 -17976
rect 3150 -18846 3160 -17976
rect 3286 -18846 3296 -17976
rect 3468 -18846 3478 -17976
rect 3604 -18846 3614 -17976
rect 3782 -18846 3792 -17976
rect 3918 -18846 3928 -17976
rect 3966 -18164 4116 -18152
rect 3962 -18648 3972 -18164
rect 4110 -18648 4120 -18164
rect 3966 -18660 4116 -18648
rect 4160 -18844 4170 -17974
rect 4296 -18844 4306 -17974
rect 4478 -18844 4488 -17974
rect 4614 -18844 4624 -17974
rect 4792 -18846 4802 -17976
rect 4928 -18846 4938 -17976
rect 5108 -18846 5118 -17976
rect 5244 -18846 5254 -17976
rect 5426 -18846 5436 -17976
rect 5562 -18846 5572 -17976
rect 5740 -18846 5750 -17976
rect 5876 -18846 5886 -17976
rect -3923 -19074 5782 -18920
rect -3552 -20060 -3542 -19190
rect -3416 -20060 -3406 -19190
rect -3234 -20060 -3224 -19190
rect -3098 -20060 -3088 -19190
rect -2920 -20062 -2910 -19192
rect -2784 -20062 -2774 -19192
rect -2604 -20062 -2594 -19192
rect -2468 -20062 -2458 -19192
rect -2286 -20062 -2276 -19192
rect -2150 -20062 -2140 -19192
rect -1566 -20060 -1556 -19190
rect -1430 -20060 -1420 -19190
rect -1248 -20060 -1238 -19190
rect -1112 -20060 -1102 -19190
rect -934 -20062 -924 -19192
rect -798 -20062 -788 -19192
rect -618 -20062 -608 -19192
rect -482 -20062 -472 -19192
rect -300 -20062 -290 -19192
rect -164 -20062 -154 -19192
rect 396 -20060 406 -19190
rect 532 -20060 542 -19190
rect 714 -20060 724 -19190
rect 850 -20060 860 -19190
rect 1028 -20062 1038 -19192
rect 1164 -20062 1174 -19192
rect 1344 -20062 1354 -19192
rect 1480 -20062 1490 -19192
rect 1662 -20062 1672 -19192
rect 1798 -20062 1808 -19192
rect 2358 -20066 2368 -19196
rect 2494 -20066 2504 -19196
rect 2676 -20066 2686 -19196
rect 2812 -20066 2822 -19196
rect 2990 -20068 3000 -19198
rect 3126 -20068 3136 -19198
rect 3306 -20068 3316 -19198
rect 3442 -20068 3452 -19198
rect 3624 -20068 3634 -19198
rect 3760 -20068 3770 -19198
rect 4316 -20066 4326 -19196
rect 4452 -20066 4462 -19196
rect 4634 -20066 4644 -19196
rect 4770 -20066 4780 -19196
rect 4948 -20068 4958 -19198
rect 5084 -20068 5094 -19198
rect 5264 -20068 5274 -19198
rect 5400 -20068 5410 -19198
rect 5582 -20068 5592 -19198
rect 5718 -20068 5728 -19198
rect -3706 -21048 -3696 -20178
rect -3570 -21048 -3560 -20178
rect -3388 -21048 -3378 -20178
rect -3252 -21048 -3242 -20178
rect -3074 -21050 -3064 -20180
rect -2938 -21050 -2928 -20180
rect -2758 -21050 -2748 -20180
rect -2622 -21050 -2612 -20180
rect -2440 -21050 -2430 -20180
rect -2304 -21050 -2294 -20180
rect -2126 -21050 -2116 -20180
rect -1990 -21050 -1980 -20180
rect -1924 -20390 -1774 -20378
rect -1928 -20874 -1918 -20390
rect -1780 -20874 -1770 -20390
rect -1924 -20886 -1774 -20874
rect -1720 -21048 -1710 -20178
rect -1584 -21048 -1574 -20178
rect -1402 -21048 -1392 -20178
rect -1266 -21048 -1256 -20178
rect -1088 -21050 -1078 -20180
rect -952 -21050 -942 -20180
rect -772 -21050 -762 -20180
rect -636 -21050 -626 -20180
rect -454 -21050 -444 -20180
rect -318 -21050 -308 -20180
rect -140 -21050 -130 -20180
rect -4 -21050 6 -20180
rect 242 -21048 252 -20178
rect 378 -21048 388 -20178
rect 560 -21048 570 -20178
rect 696 -21048 706 -20178
rect 874 -21050 884 -20180
rect 1010 -21050 1020 -20180
rect 1190 -21050 1200 -20180
rect 1326 -21050 1336 -20180
rect 1508 -21050 1518 -20180
rect 1644 -21050 1654 -20180
rect 1822 -21050 1832 -20180
rect 1958 -21050 1968 -20180
rect 2010 -20388 2160 -20376
rect 2006 -20872 2016 -20388
rect 2154 -20872 2164 -20388
rect 2010 -20884 2160 -20872
rect 2204 -21054 2214 -20184
rect 2340 -21054 2350 -20184
rect 2522 -21054 2532 -20184
rect 2658 -21054 2668 -20184
rect 2836 -21056 2846 -20186
rect 2972 -21056 2982 -20186
rect 3152 -21056 3162 -20186
rect 3288 -21056 3298 -20186
rect 3470 -21056 3480 -20186
rect 3606 -21056 3616 -20186
rect 3784 -21056 3794 -20186
rect 3920 -21056 3930 -20186
rect 4162 -21054 4172 -20184
rect 4298 -21054 4308 -20184
rect 4480 -21054 4490 -20184
rect 4616 -21054 4626 -20184
rect 4794 -21056 4804 -20186
rect 4930 -21056 4940 -20186
rect 5110 -21056 5120 -20186
rect 5246 -21056 5256 -20186
rect 5428 -21056 5438 -20186
rect 5564 -21056 5574 -20186
rect 5742 -21056 5752 -20186
rect 5878 -21056 5888 -20186
<< via1 >>
rect -5698 -7798 -5638 -7668
rect -5386 -7796 -5326 -7666
rect -5066 -7798 -5006 -7668
rect -4752 -7796 -4692 -7666
rect -4436 -7798 -4376 -7668
rect -4120 -7798 -4060 -7668
rect -3544 -8536 -3418 -7666
rect -3226 -8536 -3100 -7666
rect -2912 -8538 -2786 -7668
rect -2596 -8538 -2470 -7668
rect -2278 -8538 -2152 -7668
rect -1558 -8536 -1432 -7666
rect -1240 -8536 -1114 -7666
rect -926 -8538 -800 -7668
rect -610 -8538 -484 -7668
rect -292 -8538 -166 -7668
rect 404 -8536 530 -7666
rect 722 -8536 848 -7666
rect 1036 -8538 1162 -7668
rect 1352 -8538 1478 -7668
rect 1670 -8538 1796 -7668
rect 2366 -8542 2492 -7672
rect 2684 -8542 2810 -7672
rect 2998 -8544 3124 -7674
rect 3314 -8544 3440 -7674
rect 3632 -8544 3758 -7674
rect 4324 -8542 4450 -7672
rect 4642 -8542 4768 -7672
rect 4956 -8544 5082 -7674
rect 5272 -8544 5398 -7674
rect 5590 -8544 5716 -7674
rect -5544 -9500 -5484 -9370
rect -5226 -9500 -5166 -9370
rect -4910 -9500 -4850 -9370
rect -4598 -9502 -4538 -9372
rect -4282 -9502 -4222 -9372
rect -3698 -9524 -3572 -8654
rect -3380 -9524 -3254 -8654
rect -3066 -9526 -2940 -8656
rect -2750 -9526 -2624 -8656
rect -2432 -9526 -2306 -8656
rect -2118 -9526 -1992 -8656
rect -1712 -9524 -1586 -8654
rect -1394 -9524 -1268 -8654
rect -1080 -9526 -954 -8656
rect -764 -9526 -638 -8656
rect -446 -9526 -320 -8656
rect -132 -9526 -6 -8656
rect 60 -9370 198 -8886
rect 250 -9524 376 -8654
rect 568 -9524 694 -8654
rect 882 -9526 1008 -8656
rect 1198 -9526 1324 -8656
rect 1516 -9526 1642 -8656
rect 1830 -9526 1956 -8656
rect 2212 -9530 2338 -8660
rect 2530 -9530 2656 -8660
rect 2844 -9532 2970 -8662
rect 3160 -9532 3286 -8662
rect 3478 -9532 3604 -8662
rect 3792 -9532 3918 -8662
rect 3972 -9362 4110 -8878
rect 4170 -9530 4296 -8660
rect 4488 -9530 4614 -8660
rect 4802 -9532 4928 -8662
rect 5118 -9532 5244 -8662
rect 5436 -9532 5562 -8662
rect 5750 -9532 5876 -8662
rect -5542 -10038 -5482 -9908
rect -5226 -10036 -5166 -9906
rect -4912 -10036 -4852 -9906
rect -4596 -10034 -4536 -9904
rect -4282 -10034 -4222 -9904
rect -3916 -9948 -3776 -9626
rect -5702 -11678 -5642 -11548
rect -5386 -11676 -5326 -11546
rect -5072 -11678 -5012 -11548
rect -4752 -11680 -4692 -11550
rect -4436 -11680 -4376 -11550
rect -4120 -11680 -4060 -11550
rect -5448 -12580 -5388 -12450
rect -5136 -12580 -5076 -12450
rect -4754 -12572 -4694 -12442
rect -4436 -12578 -4376 -12448
rect -4124 -12578 -4064 -12448
rect -5292 -13056 -5232 -12926
rect -5896 -15120 -5756 -14916
rect -5454 -13800 -5394 -13670
rect -5292 -13798 -5232 -13668
rect -5136 -13802 -5076 -13672
rect -3544 -10772 -3418 -9902
rect -3226 -10772 -3100 -9902
rect -2912 -10774 -2786 -9904
rect -2596 -10774 -2470 -9904
rect -2278 -10774 -2152 -9904
rect -1558 -10772 -1432 -9902
rect -1240 -10772 -1114 -9902
rect -926 -10774 -800 -9904
rect -610 -10774 -484 -9904
rect -292 -10774 -166 -9904
rect 404 -10772 530 -9902
rect 722 -10772 848 -9902
rect 1036 -10774 1162 -9904
rect 1352 -10774 1478 -9904
rect 1670 -10774 1796 -9904
rect 2366 -10778 2492 -9908
rect 2684 -10778 2810 -9908
rect 2998 -10780 3124 -9910
rect 3314 -10780 3440 -9910
rect 3632 -10780 3758 -9910
rect 4324 -10778 4450 -9908
rect 4642 -10778 4768 -9908
rect 4956 -10780 5082 -9910
rect 5272 -10780 5398 -9910
rect 5590 -10780 5716 -9910
rect -3698 -11760 -3572 -10890
rect -3380 -11760 -3254 -10890
rect -3066 -11762 -2940 -10892
rect -2750 -11762 -2624 -10892
rect -2432 -11762 -2306 -10892
rect -2118 -11762 -1992 -10892
rect -1920 -11598 -1782 -11114
rect -1712 -11760 -1586 -10890
rect -1394 -11760 -1268 -10890
rect -1080 -11762 -954 -10892
rect -764 -11762 -638 -10892
rect -446 -11762 -320 -10892
rect -132 -11762 -6 -10892
rect 250 -11760 376 -10890
rect 568 -11760 694 -10890
rect 882 -11762 1008 -10892
rect 1198 -11762 1324 -10892
rect 1516 -11762 1642 -10892
rect 1830 -11762 1956 -10892
rect 2016 -11598 2154 -11114
rect 2212 -11766 2338 -10896
rect 2530 -11766 2656 -10896
rect 2844 -11768 2970 -10898
rect 3160 -11768 3286 -10898
rect 3478 -11768 3604 -10898
rect 3792 -11768 3918 -10898
rect 4170 -11766 4296 -10896
rect 4488 -11766 4614 -10896
rect 4802 -11768 4928 -10898
rect 5118 -11768 5244 -10898
rect 5436 -11768 5562 -10898
rect 5750 -11768 5876 -10898
rect -3544 -13008 -3418 -12138
rect -3226 -13008 -3100 -12138
rect -2912 -13010 -2786 -12140
rect -2596 -13010 -2470 -12140
rect -2278 -13010 -2152 -12140
rect -1558 -13008 -1432 -12138
rect -1240 -13008 -1114 -12138
rect -926 -13010 -800 -12140
rect -610 -13010 -484 -12140
rect -292 -13010 -166 -12140
rect 404 -13008 530 -12138
rect 722 -13008 848 -12138
rect 1036 -13010 1162 -12140
rect 1352 -13010 1478 -12140
rect 1670 -13010 1796 -12140
rect 2366 -13014 2492 -12144
rect 2684 -13014 2810 -12144
rect 2998 -13016 3124 -12146
rect 3314 -13016 3440 -12146
rect 3632 -13016 3758 -12146
rect 4324 -13014 4450 -12144
rect 4642 -13014 4768 -12144
rect 4956 -13016 5082 -12146
rect 5272 -13016 5398 -12146
rect 5590 -13016 5716 -12146
rect -3698 -13996 -3572 -13126
rect -3380 -13996 -3254 -13126
rect -3066 -13998 -2940 -13128
rect -2750 -13998 -2624 -13128
rect -2432 -13998 -2306 -13128
rect -2118 -13998 -1992 -13128
rect -1712 -13996 -1586 -13126
rect -1394 -13996 -1268 -13126
rect -1080 -13998 -954 -13128
rect -764 -13998 -638 -13128
rect -446 -13998 -320 -13128
rect -132 -13998 -6 -13128
rect 58 -13848 196 -13364
rect 250 -13996 376 -13126
rect 568 -13996 694 -13126
rect 882 -13998 1008 -13128
rect 1198 -13998 1324 -13128
rect 1516 -13998 1642 -13128
rect 1830 -13998 1956 -13128
rect 2212 -14002 2338 -13132
rect 2530 -14002 2656 -13132
rect 2844 -14004 2970 -13134
rect 3160 -14004 3286 -13134
rect 3478 -14004 3604 -13134
rect 3792 -14004 3918 -13134
rect 3974 -13852 4112 -13368
rect 4170 -14002 4296 -13132
rect 4488 -14002 4614 -13132
rect 4802 -14004 4928 -13134
rect 5118 -14004 5244 -13134
rect 5436 -14004 5562 -13134
rect 5750 -14004 5876 -13134
rect -4594 -14248 -4534 -14118
rect -4274 -14246 -4214 -14116
rect -4646 -14662 -4538 -14540
rect -4271 -15007 -4197 -14933
rect -4694 -15624 -4634 -15494
rect -4376 -15624 -4316 -15494
rect -5400 -16318 -5330 -16184
rect -4850 -16316 -4790 -16186
rect -4530 -16314 -4470 -16184
rect -4220 -16320 -4160 -16190
rect -3544 -15244 -3418 -14374
rect -3226 -15244 -3100 -14374
rect -2912 -15246 -2786 -14376
rect -2596 -15246 -2470 -14376
rect -2278 -15246 -2152 -14376
rect -1558 -15244 -1432 -14374
rect -1240 -15244 -1114 -14374
rect -926 -15246 -800 -14376
rect -610 -15246 -484 -14376
rect -292 -15246 -166 -14376
rect 404 -15244 530 -14374
rect 722 -15244 848 -14374
rect 1036 -15246 1162 -14376
rect 1352 -15246 1478 -14376
rect 1670 -15246 1796 -14376
rect 2366 -15250 2492 -14380
rect 2684 -15250 2810 -14380
rect 2998 -15252 3124 -14382
rect 3314 -15252 3440 -14382
rect 3632 -15252 3758 -14382
rect 4324 -15250 4450 -14380
rect 4642 -15250 4768 -14380
rect 4956 -15252 5082 -14382
rect 5272 -15252 5398 -14382
rect 5590 -15252 5716 -14382
rect -3698 -16232 -3572 -15362
rect -3380 -16232 -3254 -15362
rect -3066 -16234 -2940 -15364
rect -2750 -16234 -2624 -15364
rect -2432 -16234 -2306 -15364
rect -2118 -16234 -1992 -15364
rect -1924 -16036 -1786 -15552
rect -1712 -16232 -1586 -15362
rect -1394 -16232 -1268 -15362
rect -1080 -16234 -954 -15364
rect -764 -16234 -638 -15364
rect -446 -16234 -320 -15364
rect -132 -16234 -6 -15364
rect 250 -16232 376 -15362
rect 568 -16232 694 -15362
rect 882 -16234 1008 -15364
rect 1198 -16234 1324 -15364
rect 1516 -16234 1642 -15364
rect 1830 -16234 1956 -15364
rect 2022 -16044 2160 -15560
rect 2212 -16238 2338 -15368
rect 2530 -16238 2656 -15368
rect 2844 -16240 2970 -15370
rect 3160 -16240 3286 -15370
rect 3478 -16240 3604 -15370
rect 3792 -16240 3918 -15370
rect 4170 -16238 4296 -15368
rect 4488 -16238 4614 -15368
rect 4802 -16240 4928 -15370
rect 5118 -16240 5244 -15370
rect 5436 -16240 5562 -15370
rect 5750 -16240 5876 -15370
rect -5542 -17124 -5482 -16994
rect -5228 -17124 -5168 -16994
rect -4912 -17126 -4852 -16996
rect -4594 -17126 -4534 -16996
rect -4276 -17128 -4216 -16998
rect -3908 -17170 -3786 -16912
rect -5702 -18774 -5642 -18644
rect -5386 -18776 -5326 -18646
rect -5068 -18776 -5008 -18646
rect -4752 -18776 -4692 -18646
rect -4436 -18776 -4376 -18646
rect -4118 -18776 -4058 -18646
rect -3544 -17850 -3418 -16980
rect -3226 -17850 -3100 -16980
rect -2912 -17852 -2786 -16982
rect -2596 -17852 -2470 -16982
rect -2278 -17852 -2152 -16982
rect -1558 -17850 -1432 -16980
rect -1240 -17850 -1114 -16980
rect -926 -17852 -800 -16982
rect -610 -17852 -484 -16982
rect -292 -17852 -166 -16982
rect 404 -17850 530 -16980
rect 722 -17850 848 -16980
rect 1036 -17852 1162 -16982
rect 1352 -17852 1478 -16982
rect 1670 -17852 1796 -16982
rect 2366 -17856 2492 -16986
rect 2684 -17856 2810 -16986
rect 2998 -17858 3124 -16988
rect 3314 -17858 3440 -16988
rect 3632 -17858 3758 -16988
rect 4324 -17856 4450 -16986
rect 4642 -17856 4768 -16986
rect 4956 -17858 5082 -16988
rect 5272 -17858 5398 -16988
rect 5590 -17858 5716 -16988
rect -3698 -18838 -3572 -17968
rect -3380 -18838 -3254 -17968
rect -3066 -18840 -2940 -17970
rect -2750 -18840 -2624 -17970
rect -2432 -18840 -2306 -17970
rect -2118 -18840 -1992 -17970
rect -1712 -18838 -1586 -17968
rect -1394 -18838 -1268 -17968
rect -1080 -18840 -954 -17970
rect -764 -18840 -638 -17970
rect -446 -18840 -320 -17970
rect -132 -18840 -6 -17970
rect 56 -18648 194 -18164
rect 250 -18838 376 -17968
rect 568 -18838 694 -17968
rect 882 -18840 1008 -17970
rect 1198 -18840 1324 -17970
rect 1516 -18840 1642 -17970
rect 1830 -18840 1956 -17970
rect 2212 -18844 2338 -17974
rect 2530 -18844 2656 -17974
rect 2844 -18846 2970 -17976
rect 3160 -18846 3286 -17976
rect 3478 -18846 3604 -17976
rect 3792 -18846 3918 -17976
rect 3972 -18648 4110 -18164
rect 4170 -18844 4296 -17974
rect 4488 -18844 4614 -17974
rect 4802 -18846 4928 -17976
rect 5118 -18846 5244 -17976
rect 5436 -18846 5562 -17976
rect 5750 -18846 5876 -17976
rect -3542 -20060 -3416 -19190
rect -3224 -20060 -3098 -19190
rect -2910 -20062 -2784 -19192
rect -2594 -20062 -2468 -19192
rect -2276 -20062 -2150 -19192
rect -1556 -20060 -1430 -19190
rect -1238 -20060 -1112 -19190
rect -924 -20062 -798 -19192
rect -608 -20062 -482 -19192
rect -290 -20062 -164 -19192
rect 406 -20060 532 -19190
rect 724 -20060 850 -19190
rect 1038 -20062 1164 -19192
rect 1354 -20062 1480 -19192
rect 1672 -20062 1798 -19192
rect 2368 -20066 2494 -19196
rect 2686 -20066 2812 -19196
rect 3000 -20068 3126 -19198
rect 3316 -20068 3442 -19198
rect 3634 -20068 3760 -19198
rect 4326 -20066 4452 -19196
rect 4644 -20066 4770 -19196
rect 4958 -20068 5084 -19198
rect 5274 -20068 5400 -19198
rect 5592 -20068 5718 -19198
rect -3696 -21048 -3570 -20178
rect -3378 -21048 -3252 -20178
rect -3064 -21050 -2938 -20180
rect -2748 -21050 -2622 -20180
rect -2430 -21050 -2304 -20180
rect -2116 -21050 -1990 -20180
rect -1918 -20874 -1780 -20390
rect -1710 -21048 -1584 -20178
rect -1392 -21048 -1266 -20178
rect -1078 -21050 -952 -20180
rect -762 -21050 -636 -20180
rect -444 -21050 -318 -20180
rect -130 -21050 -4 -20180
rect 252 -21048 378 -20178
rect 570 -21048 696 -20178
rect 884 -21050 1010 -20180
rect 1200 -21050 1326 -20180
rect 1518 -21050 1644 -20180
rect 1832 -21050 1958 -20180
rect 2016 -20872 2154 -20388
rect 2214 -21054 2340 -20184
rect 2532 -21054 2658 -20184
rect 2846 -21056 2972 -20186
rect 3162 -21056 3288 -20186
rect 3480 -21056 3606 -20186
rect 3794 -21056 3920 -20186
rect 4172 -21054 4298 -20184
rect 4490 -21054 4616 -20184
rect 4804 -21056 4930 -20186
rect 5120 -21056 5246 -20186
rect 5438 -21056 5564 -20186
rect 5752 -21056 5878 -20186
<< metal2 >>
rect -5698 -7668 -5638 -7658
rect -5386 -7666 -5326 -7656
rect -5638 -7770 -5386 -7690
rect -5698 -7808 -5638 -7798
rect -5066 -7668 -5006 -7658
rect -5326 -7770 -5066 -7690
rect -5386 -7806 -5326 -7796
rect -4752 -7666 -4692 -7656
rect -5006 -7770 -4752 -7690
rect -5066 -7808 -5006 -7798
rect -4436 -7668 -4376 -7658
rect -4692 -7770 -4436 -7690
rect -4752 -7806 -4692 -7796
rect -4120 -7668 -4060 -7658
rect -4376 -7770 -4120 -7692
rect -4436 -7808 -4376 -7798
rect -3544 -7666 -3418 -7656
rect -4060 -7770 -3825 -7692
rect -4120 -7808 -4060 -7798
rect -3903 -8667 -3825 -7770
rect -3226 -7666 -3100 -7656
rect -3418 -8362 -3226 -7828
rect -3544 -8546 -3418 -8536
rect -2912 -7668 -2786 -7658
rect -3100 -8362 -2912 -7828
rect -3226 -8546 -3100 -8536
rect -2596 -7668 -2470 -7658
rect -2786 -8362 -2596 -7828
rect -2912 -8548 -2786 -8538
rect -2278 -7668 -2152 -7658
rect -2470 -8362 -2278 -7828
rect -2596 -8548 -2470 -8538
rect -1558 -7666 -1432 -7656
rect -2152 -8362 -1558 -7828
rect -2278 -8548 -2152 -8538
rect -1240 -7666 -1114 -7656
rect -1432 -8362 -1240 -7828
rect -1558 -8546 -1432 -8536
rect -926 -7668 -800 -7658
rect -1114 -8362 -926 -7828
rect -1240 -8546 -1114 -8536
rect -610 -7668 -484 -7658
rect -800 -8362 -610 -7828
rect -926 -8548 -800 -8538
rect -292 -7668 -166 -7658
rect -484 -8362 -292 -7828
rect -610 -8548 -484 -8538
rect 404 -7666 530 -7656
rect -166 -8362 404 -7828
rect -292 -8548 -166 -8538
rect 722 -7666 848 -7656
rect 530 -8362 722 -7828
rect 404 -8546 530 -8536
rect 1036 -7668 1162 -7658
rect 848 -8362 1036 -7828
rect 722 -8546 848 -8536
rect 1352 -7668 1478 -7658
rect 1162 -8362 1352 -7828
rect 1036 -8548 1162 -8538
rect 1670 -7668 1796 -7658
rect 1478 -8362 1670 -7828
rect 1352 -8548 1478 -8538
rect 2366 -7672 2492 -7662
rect 1796 -8362 2366 -7828
rect 1670 -8548 1796 -8538
rect 2684 -7672 2810 -7662
rect 2492 -8362 2684 -7828
rect 2366 -8552 2492 -8542
rect 2998 -7674 3124 -7664
rect 2810 -8362 2998 -7828
rect 2684 -8552 2810 -8542
rect 3314 -7674 3440 -7664
rect 3124 -8362 3314 -7828
rect 2998 -8554 3124 -8544
rect 3632 -7674 3758 -7664
rect 3440 -8362 3632 -7828
rect 3314 -8554 3440 -8544
rect 4324 -7672 4450 -7662
rect 3758 -7846 4324 -7828
rect 4642 -7672 4768 -7662
rect 4450 -7846 4642 -7828
rect 4956 -7674 5082 -7664
rect 4768 -7846 4956 -7828
rect 5272 -7674 5398 -7664
rect 5082 -7846 5272 -7828
rect 5590 -7674 5716 -7664
rect 5398 -7846 5590 -7828
rect 3758 -8356 3808 -7846
rect 3758 -8362 4324 -8356
rect 3808 -8366 4324 -8362
rect 3632 -8554 3758 -8544
rect 4450 -8366 4642 -8356
rect 4324 -8552 4450 -8542
rect 4768 -8366 4956 -8356
rect 4642 -8552 4768 -8542
rect 5082 -8366 5272 -8356
rect 4956 -8554 5082 -8544
rect 5398 -8366 5590 -8356
rect 5272 -8554 5398 -8544
rect 5590 -8554 5716 -8544
rect -3698 -8654 -3572 -8644
rect -3903 -8745 -3698 -8667
rect -5544 -9370 -5484 -9360
rect -5226 -9370 -5166 -9360
rect -5484 -9478 -5226 -9394
rect -5544 -9510 -5484 -9500
rect -4910 -9370 -4850 -9360
rect -5166 -9478 -4910 -9394
rect -5226 -9510 -5166 -9500
rect -4598 -9372 -4538 -9362
rect -4850 -9478 -4598 -9394
rect -4910 -9510 -4850 -9500
rect -4282 -9372 -4222 -9362
rect -4538 -9478 -4282 -9394
rect -4598 -9512 -4538 -9502
rect -4222 -9478 -3848 -9394
rect -4282 -9512 -4222 -9502
rect -3932 -9616 -3848 -9478
rect -3380 -8654 -3254 -8644
rect -3572 -9374 -3380 -8888
rect -3698 -9534 -3572 -9524
rect -3066 -8656 -2940 -8646
rect -3254 -9022 -3066 -8888
rect -2750 -8656 -2624 -8646
rect -2940 -9022 -2750 -8888
rect -2432 -8656 -2306 -8646
rect -2624 -9022 -2432 -8888
rect -2118 -8656 -1992 -8646
rect -2306 -9022 -2118 -8888
rect -1712 -8654 -1586 -8644
rect -1992 -9022 -1712 -8888
rect -1394 -8654 -1268 -8644
rect -1586 -9022 -1394 -8888
rect -1080 -8656 -954 -8646
rect -1268 -9022 -1080 -8888
rect -764 -8656 -638 -8646
rect -954 -9022 -764 -8888
rect -446 -8656 -320 -8646
rect -638 -9022 -446 -8888
rect -132 -8656 -6 -8646
rect -320 -9022 -132 -8888
rect -3254 -9336 -3202 -9022
rect -3254 -9374 -3066 -9336
rect -3380 -9534 -3254 -9524
rect -2940 -9374 -2750 -9336
rect -3066 -9536 -2940 -9526
rect -2624 -9374 -2432 -9336
rect -2750 -9536 -2624 -9526
rect -2306 -9374 -2118 -9336
rect -2432 -9536 -2306 -9526
rect -1992 -9374 -1712 -9336
rect -2118 -9536 -1992 -9526
rect -1586 -9374 -1394 -9336
rect -1712 -9534 -1586 -9524
rect -1268 -9374 -1080 -9336
rect -1394 -9534 -1268 -9524
rect -954 -9374 -764 -9336
rect -1080 -9536 -954 -9526
rect -638 -9374 -446 -9336
rect -764 -9536 -638 -9526
rect -320 -9374 -132 -9336
rect -446 -9536 -320 -9526
rect 250 -8654 376 -8644
rect 60 -8886 198 -8876
rect -6 -9022 60 -8888
rect -6 -9370 60 -9336
rect 198 -9022 250 -8888
rect 198 -9370 250 -9336
rect -6 -9374 250 -9370
rect 60 -9380 198 -9374
rect -132 -9536 -6 -9526
rect 568 -8654 694 -8644
rect 376 -9022 568 -8888
rect 376 -9374 568 -9336
rect 250 -9534 376 -9524
rect 882 -8656 1008 -8646
rect 694 -9022 882 -8888
rect 694 -9374 882 -9336
rect 568 -9534 694 -9524
rect 1198 -8656 1324 -8646
rect 1008 -9022 1198 -8888
rect 1008 -9374 1198 -9336
rect 882 -9536 1008 -9526
rect 1516 -8656 1642 -8646
rect 1324 -9022 1516 -8888
rect 1324 -9374 1516 -9336
rect 1198 -9536 1324 -9526
rect 1830 -8656 1956 -8646
rect 1642 -9022 1830 -8888
rect 1642 -9374 1830 -9336
rect 1516 -9536 1642 -9526
rect 2212 -8660 2338 -8650
rect 1956 -9022 2212 -8888
rect 1956 -9374 2212 -9336
rect 1830 -9536 1956 -9526
rect 2530 -8660 2656 -8650
rect 2338 -9022 2530 -8888
rect 2338 -9374 2530 -9336
rect 2212 -9540 2338 -9530
rect 2844 -8662 2970 -8652
rect 2656 -9022 2844 -8888
rect 2656 -9374 2844 -9336
rect 2530 -9540 2656 -9530
rect 3160 -8662 3286 -8652
rect 2970 -9022 3160 -8888
rect 2970 -9374 3160 -9336
rect 2844 -9542 2970 -9532
rect 3478 -8662 3604 -8652
rect 3286 -9022 3478 -8888
rect 3332 -9336 3478 -9022
rect 3286 -9374 3478 -9336
rect 3160 -9542 3286 -9532
rect 3792 -8662 3918 -8652
rect 3604 -9374 3792 -8888
rect 3478 -9542 3604 -9532
rect 4170 -8660 4296 -8650
rect 3972 -8878 4110 -8868
rect 3918 -9362 3972 -8888
rect 4110 -9362 4170 -8888
rect 3918 -9374 4170 -9362
rect 3792 -9542 3918 -9532
rect 4488 -8660 4614 -8650
rect 4296 -9374 4488 -8888
rect 4170 -9540 4296 -9530
rect 4802 -8662 4928 -8652
rect 4614 -9374 4802 -8888
rect 4488 -9540 4614 -9530
rect 5118 -8662 5244 -8652
rect 4928 -9374 5118 -8888
rect 4802 -9542 4928 -9532
rect 5436 -8662 5562 -8652
rect 5244 -9374 5436 -8888
rect 5118 -9542 5244 -9532
rect 5750 -8662 5876 -8652
rect 5562 -9374 5750 -8888
rect 5436 -9542 5562 -9532
rect 5750 -9542 5876 -9532
rect -3932 -9626 -3776 -9616
rect -5542 -9908 -5482 -9898
rect -5226 -9906 -5166 -9896
rect -5482 -10008 -5226 -9924
rect -5542 -10048 -5482 -10038
rect -4912 -9906 -4852 -9896
rect -5166 -10008 -4912 -9924
rect -5226 -10046 -5166 -10036
rect -4596 -9904 -4536 -9894
rect -4852 -10008 -4596 -9924
rect -4912 -10046 -4852 -10036
rect -4282 -9904 -4222 -9894
rect -4536 -10008 -4282 -9924
rect -4596 -10044 -4536 -10034
rect -3932 -9924 -3916 -9626
rect -4222 -9948 -3916 -9924
rect -4222 -9958 -3776 -9948
rect -3544 -9902 -3418 -9892
rect -4222 -10008 -3848 -9958
rect -4282 -10044 -4222 -10034
rect -3226 -9902 -3100 -9892
rect -3418 -10614 -3226 -10080
rect -3544 -10782 -3418 -10772
rect -2912 -9904 -2786 -9894
rect -3100 -10614 -2912 -10080
rect -3226 -10782 -3100 -10772
rect -2596 -9904 -2470 -9894
rect -2786 -10614 -2596 -10080
rect -2912 -10784 -2786 -10774
rect -2278 -9904 -2152 -9894
rect -2470 -10614 -2278 -10080
rect -2596 -10784 -2470 -10774
rect -1558 -9902 -1432 -9892
rect -2152 -10614 -1558 -10080
rect -2278 -10784 -2152 -10774
rect -1240 -9902 -1114 -9892
rect -1432 -10614 -1240 -10080
rect -1558 -10782 -1432 -10772
rect -926 -9904 -800 -9894
rect -1114 -10614 -926 -10080
rect -1240 -10782 -1114 -10772
rect -610 -9904 -484 -9894
rect -800 -10614 -610 -10080
rect -926 -10784 -800 -10774
rect -292 -9904 -166 -9894
rect -484 -10614 -292 -10080
rect -610 -10784 -484 -10774
rect 404 -9902 530 -9892
rect -166 -10614 404 -10080
rect -292 -10784 -166 -10774
rect 722 -9902 848 -9892
rect 530 -10614 722 -10080
rect 404 -10782 530 -10772
rect 1036 -9904 1162 -9894
rect 848 -10614 1036 -10080
rect 722 -10782 848 -10772
rect 1352 -9904 1478 -9894
rect 1162 -10614 1352 -10080
rect 1036 -10784 1162 -10774
rect 1670 -9904 1796 -9894
rect 1478 -10614 1670 -10080
rect 1352 -10784 1478 -10774
rect 2366 -9908 2492 -9898
rect 1796 -10614 2366 -10080
rect 1670 -10784 1796 -10774
rect 2684 -9908 2810 -9898
rect 2492 -10614 2684 -10080
rect 2366 -10788 2492 -10778
rect 2998 -9910 3124 -9900
rect 2810 -10614 2998 -10080
rect 2684 -10788 2810 -10778
rect 3314 -9910 3440 -9900
rect 3124 -10614 3314 -10080
rect 2998 -10790 3124 -10780
rect 3632 -9910 3758 -9900
rect 3440 -10614 3632 -10080
rect 3314 -10790 3440 -10780
rect 4324 -9908 4450 -9898
rect 3758 -10092 4324 -10080
rect 4642 -9908 4768 -9898
rect 4450 -10092 4642 -10080
rect 4956 -9910 5082 -9900
rect 4768 -10092 4956 -10080
rect 5272 -9910 5398 -9900
rect 5082 -10092 5272 -10080
rect 5590 -9910 5716 -9900
rect 5398 -10092 5590 -10080
rect 3758 -10602 3808 -10092
rect 3758 -10614 4324 -10602
rect 3632 -10790 3758 -10780
rect 4450 -10614 4642 -10602
rect 4324 -10788 4450 -10778
rect 4768 -10614 4956 -10602
rect 4642 -10788 4768 -10778
rect 5082 -10614 5272 -10602
rect 4956 -10790 5082 -10780
rect 5398 -10614 5590 -10602
rect 5272 -10790 5398 -10780
rect 5590 -10790 5716 -10780
rect -3890 -10890 -3730 -10888
rect -3698 -10890 -3572 -10880
rect -5702 -11548 -5642 -11538
rect -5386 -11546 -5326 -11536
rect -5642 -11656 -5386 -11572
rect -5702 -11688 -5642 -11678
rect -5072 -11548 -5012 -11538
rect -5326 -11656 -5072 -11572
rect -5386 -11686 -5326 -11676
rect -4752 -11550 -4692 -11540
rect -5012 -11656 -4752 -11572
rect -5072 -11688 -5012 -11678
rect -4436 -11550 -4376 -11540
rect -4692 -11656 -4436 -11572
rect -4752 -11690 -4692 -11680
rect -4120 -11550 -4060 -11540
rect -4376 -11656 -4120 -11572
rect -4436 -11690 -4376 -11680
rect -3890 -11572 -3698 -10890
rect -4060 -11656 -3698 -11572
rect -4120 -11690 -4060 -11680
rect -3889 -11760 -3698 -11656
rect -3380 -10890 -3254 -10880
rect -3572 -11600 -3380 -11114
rect -3889 -11770 -3572 -11760
rect -3066 -10892 -2940 -10882
rect -3254 -11234 -3066 -11114
rect -2750 -10892 -2624 -10882
rect -2940 -11234 -2750 -11114
rect -2432 -10892 -2306 -10882
rect -2624 -11234 -2432 -11114
rect -2118 -10892 -1992 -10882
rect -2306 -11234 -2118 -11114
rect -1712 -10890 -1586 -10880
rect -1920 -11114 -1782 -11104
rect -1992 -11234 -1920 -11114
rect -1782 -11234 -1712 -11114
rect -1394 -10890 -1268 -10880
rect -1586 -11234 -1394 -11114
rect -1080 -10892 -954 -10882
rect -1268 -11234 -1080 -11114
rect -764 -10892 -638 -10882
rect -954 -11234 -764 -11114
rect -446 -10892 -320 -10882
rect -638 -11234 -446 -11114
rect -132 -10892 -6 -10882
rect -320 -11234 -132 -11114
rect -3254 -11548 -3214 -11234
rect -3254 -11600 -3066 -11548
rect -3380 -11770 -3254 -11760
rect -2940 -11600 -2750 -11548
rect -3889 -11772 -3654 -11770
rect -3066 -11772 -2940 -11762
rect -2624 -11600 -2432 -11548
rect -2750 -11772 -2624 -11762
rect -2306 -11600 -2118 -11548
rect -2432 -11772 -2306 -11762
rect -1992 -11598 -1920 -11548
rect -1782 -11598 -1712 -11548
rect -1992 -11600 -1712 -11598
rect -1920 -11608 -1782 -11600
rect -2118 -11772 -1992 -11762
rect -1586 -11600 -1394 -11548
rect -1712 -11770 -1586 -11760
rect -1268 -11600 -1080 -11548
rect -1394 -11770 -1268 -11760
rect -954 -11600 -764 -11548
rect -1080 -11772 -954 -11762
rect -638 -11600 -446 -11548
rect -764 -11772 -638 -11762
rect -320 -11600 -132 -11548
rect -446 -11772 -320 -11762
rect 250 -10890 376 -10880
rect -6 -11234 250 -11114
rect -6 -11600 250 -11548
rect -132 -11772 -6 -11762
rect 568 -10890 694 -10880
rect 376 -11234 568 -11114
rect 376 -11600 568 -11548
rect 250 -11770 376 -11760
rect 882 -10892 1008 -10882
rect 694 -11234 882 -11114
rect 694 -11600 882 -11548
rect 568 -11770 694 -11760
rect 1198 -10892 1324 -10882
rect 1008 -11234 1198 -11114
rect 1008 -11600 1198 -11548
rect 882 -11772 1008 -11762
rect 1516 -10892 1642 -10882
rect 1324 -11234 1516 -11114
rect 1324 -11600 1516 -11548
rect 1198 -11772 1324 -11762
rect 1830 -10892 1956 -10882
rect 1642 -11234 1830 -11114
rect 1642 -11600 1830 -11548
rect 1516 -11772 1642 -11762
rect 2212 -10896 2338 -10886
rect 2016 -11114 2154 -11104
rect 1956 -11234 2016 -11114
rect 1956 -11598 2016 -11548
rect 2154 -11234 2212 -11114
rect 2154 -11598 2212 -11548
rect 1956 -11600 2212 -11598
rect 2016 -11608 2154 -11600
rect 1830 -11772 1956 -11762
rect 2530 -10896 2656 -10886
rect 2338 -11234 2530 -11114
rect 2338 -11600 2530 -11548
rect -5448 -12450 -5388 -12440
rect -5136 -12450 -5076 -12440
rect -5388 -12550 -5136 -12472
rect -5448 -12590 -5388 -12580
rect -4754 -12442 -4694 -12432
rect -5076 -12550 -4754 -12472
rect -5136 -12590 -5076 -12580
rect -5292 -12926 -5232 -12916
rect -5606 -13036 -5292 -12958
rect -5606 -14563 -5528 -13036
rect -5292 -13066 -5232 -13056
rect -4977 -13403 -4899 -12550
rect -4436 -12448 -4376 -12438
rect -4694 -12550 -4436 -12472
rect -4754 -12582 -4694 -12572
rect -4124 -12448 -4064 -12438
rect -4376 -12550 -4124 -12472
rect -4436 -12588 -4376 -12578
rect -3889 -12472 -3811 -11772
rect 2212 -11776 2338 -11766
rect 2844 -10898 2970 -10888
rect 2656 -11234 2844 -11114
rect 2656 -11600 2844 -11548
rect 2530 -11776 2656 -11766
rect 3160 -10898 3286 -10888
rect 2970 -11234 3160 -11114
rect 2970 -11600 3160 -11548
rect 2844 -11778 2970 -11768
rect 3478 -10898 3604 -10888
rect 3286 -11234 3478 -11114
rect 3320 -11548 3478 -11234
rect 3286 -11600 3478 -11548
rect 3160 -11778 3286 -11768
rect 3792 -10898 3918 -10888
rect 3604 -11600 3792 -11114
rect 3478 -11778 3604 -11768
rect 4170 -10896 4296 -10886
rect 3918 -11600 4170 -11114
rect 3792 -11778 3918 -11768
rect 4488 -10896 4614 -10886
rect 4296 -11600 4488 -11114
rect 4170 -11776 4296 -11766
rect 4802 -10898 4928 -10888
rect 4614 -11600 4802 -11114
rect 4488 -11776 4614 -11766
rect 5118 -10898 5244 -10888
rect 4928 -11600 5118 -11114
rect 4802 -11778 4928 -11768
rect 5436 -10898 5562 -10888
rect 5244 -11600 5436 -11114
rect 5118 -11778 5244 -11768
rect 5750 -10898 5876 -10888
rect 5562 -11600 5750 -11114
rect 5436 -11778 5562 -11768
rect 5750 -11778 5876 -11768
rect -4064 -12550 -3811 -12472
rect -3544 -12138 -3418 -12128
rect -4124 -12588 -4064 -12578
rect -3226 -12138 -3100 -12128
rect -3418 -12806 -3226 -12272
rect -3544 -13018 -3418 -13008
rect -2912 -12140 -2786 -12130
rect -3100 -12806 -2912 -12272
rect -3226 -13018 -3100 -13008
rect -2596 -12140 -2470 -12130
rect -2786 -12806 -2596 -12272
rect -2912 -13020 -2786 -13010
rect -2278 -12140 -2152 -12130
rect -2470 -12806 -2278 -12272
rect -2596 -13020 -2470 -13010
rect -1558 -12138 -1432 -12128
rect -2152 -12806 -1558 -12272
rect -2278 -13020 -2152 -13010
rect -1240 -12138 -1114 -12128
rect -1432 -12806 -1240 -12272
rect -1558 -13018 -1432 -13008
rect -926 -12140 -800 -12130
rect -1114 -12806 -926 -12272
rect -1240 -13018 -1114 -13008
rect -610 -12140 -484 -12130
rect -800 -12806 -610 -12272
rect -926 -13020 -800 -13010
rect -292 -12140 -166 -12130
rect -484 -12806 -292 -12272
rect -610 -13020 -484 -13010
rect 404 -12138 530 -12128
rect -166 -12806 404 -12272
rect -292 -13020 -166 -13010
rect 722 -12138 848 -12128
rect 530 -12806 722 -12272
rect 404 -13018 530 -13008
rect 1036 -12140 1162 -12130
rect 848 -12806 1036 -12272
rect 722 -13018 848 -13008
rect 1352 -12140 1478 -12130
rect 1162 -12806 1352 -12272
rect 1036 -13020 1162 -13010
rect 1670 -12140 1796 -12130
rect 1478 -12806 1670 -12272
rect 1352 -13020 1478 -13010
rect 2366 -12144 2492 -12134
rect 1796 -12806 2366 -12272
rect 1670 -13020 1796 -13010
rect 2684 -12144 2810 -12134
rect 2492 -12806 2684 -12272
rect 2366 -13024 2492 -13014
rect 2998 -12146 3124 -12136
rect 2810 -12806 2998 -12272
rect 2684 -13024 2810 -13014
rect 3314 -12146 3440 -12136
rect 3124 -12806 3314 -12272
rect 2998 -13026 3124 -13016
rect 3632 -12146 3758 -12136
rect 3440 -12806 3632 -12272
rect 3314 -13026 3440 -13016
rect 4324 -12144 4450 -12134
rect 3758 -12284 4324 -12272
rect 4642 -12144 4768 -12134
rect 4450 -12284 4642 -12272
rect 4956 -12146 5082 -12136
rect 4768 -12284 4956 -12272
rect 5272 -12146 5398 -12136
rect 5082 -12284 5272 -12272
rect 5590 -12146 5716 -12136
rect 5398 -12284 5590 -12272
rect 3758 -12794 3808 -12284
rect 3758 -12806 4324 -12794
rect 3632 -13026 3758 -13016
rect 4450 -12806 4642 -12794
rect 4324 -13024 4450 -13014
rect 4768 -12806 4956 -12794
rect 4642 -13024 4768 -13014
rect 5082 -12806 5272 -12794
rect 4956 -13026 5082 -13016
rect 5398 -12806 5590 -12794
rect 5272 -13026 5398 -13016
rect 5590 -13026 5716 -13016
rect -5303 -13481 -4899 -13403
rect -3698 -13126 -3572 -13116
rect -5454 -13670 -5394 -13660
rect -5454 -13810 -5394 -13800
rect -5303 -13668 -5225 -13481
rect -5303 -13798 -5292 -13668
rect -5232 -13798 -5225 -13668
rect -5303 -13815 -5225 -13798
rect -5136 -13672 -5076 -13662
rect -5136 -13812 -5076 -13802
rect -3380 -13126 -3254 -13116
rect -3572 -13852 -3380 -13366
rect -3698 -14006 -3572 -13996
rect -3066 -13128 -2940 -13118
rect -3254 -13488 -3066 -13366
rect -2750 -13128 -2624 -13118
rect -2940 -13488 -2750 -13366
rect -2432 -13128 -2306 -13118
rect -2624 -13488 -2432 -13366
rect -2118 -13128 -1992 -13118
rect -2306 -13488 -2118 -13366
rect -1712 -13126 -1586 -13116
rect -1992 -13488 -1712 -13366
rect -1394 -13126 -1268 -13116
rect -1586 -13488 -1394 -13366
rect -1080 -13128 -954 -13118
rect -1268 -13488 -1080 -13366
rect -764 -13128 -638 -13118
rect -954 -13488 -764 -13366
rect -446 -13128 -320 -13118
rect -638 -13488 -446 -13366
rect -132 -13128 -6 -13118
rect -320 -13488 -132 -13366
rect -3254 -13802 -3208 -13488
rect -3254 -13852 -3066 -13802
rect -3380 -14006 -3254 -13996
rect -2940 -13852 -2750 -13802
rect -3066 -14008 -2940 -13998
rect -2624 -13852 -2432 -13802
rect -2750 -14008 -2624 -13998
rect -2306 -13852 -2118 -13802
rect -2432 -14008 -2306 -13998
rect -1992 -13852 -1712 -13802
rect -2118 -14008 -1992 -13998
rect -1586 -13852 -1394 -13802
rect -1712 -14006 -1586 -13996
rect -1268 -13852 -1080 -13802
rect -1394 -14006 -1268 -13996
rect -954 -13852 -764 -13802
rect -1080 -14008 -954 -13998
rect -638 -13852 -446 -13802
rect -764 -14008 -638 -13998
rect -320 -13852 -132 -13802
rect -446 -14008 -320 -13998
rect 250 -13126 376 -13116
rect 58 -13364 196 -13354
rect -6 -13488 58 -13366
rect -6 -13848 58 -13802
rect 196 -13488 250 -13366
rect 196 -13848 250 -13802
rect -6 -13852 250 -13848
rect 58 -13858 196 -13852
rect -132 -14008 -6 -13998
rect 568 -13126 694 -13116
rect 376 -13488 568 -13366
rect 376 -13852 568 -13802
rect 250 -14006 376 -13996
rect 882 -13128 1008 -13118
rect 694 -13488 882 -13366
rect 694 -13852 882 -13802
rect 568 -14006 694 -13996
rect 1198 -13128 1324 -13118
rect 1008 -13488 1198 -13366
rect 1008 -13852 1198 -13802
rect 882 -14008 1008 -13998
rect 1516 -13128 1642 -13118
rect 1324 -13488 1516 -13366
rect 1324 -13852 1516 -13802
rect 1198 -14008 1324 -13998
rect 1830 -13128 1956 -13118
rect 1642 -13488 1830 -13366
rect 1642 -13852 1830 -13802
rect 1516 -14008 1642 -13998
rect 2212 -13132 2338 -13122
rect 1956 -13488 2212 -13366
rect 1956 -13852 2212 -13802
rect 1830 -14008 1956 -13998
rect 2530 -13132 2656 -13122
rect 2338 -13488 2530 -13366
rect 2338 -13852 2530 -13802
rect 2212 -14012 2338 -14002
rect 2844 -13134 2970 -13124
rect 2656 -13488 2844 -13366
rect 2656 -13852 2844 -13802
rect 2530 -14012 2656 -14002
rect 3160 -13134 3286 -13124
rect 2970 -13488 3160 -13366
rect 2970 -13852 3160 -13802
rect 2844 -14014 2970 -14004
rect 3478 -13134 3604 -13124
rect 3286 -13488 3478 -13366
rect 3326 -13802 3478 -13488
rect 3286 -13852 3478 -13802
rect 3160 -14014 3286 -14004
rect 3792 -13134 3918 -13124
rect 3604 -13852 3792 -13366
rect 3478 -14014 3604 -14004
rect 4170 -13132 4296 -13122
rect 3974 -13366 4112 -13358
rect 3918 -13368 4170 -13366
rect 3918 -13852 3974 -13368
rect 4112 -13852 4170 -13368
rect 3974 -13862 4112 -13852
rect 3792 -14014 3918 -14004
rect 4488 -13132 4614 -13122
rect 4296 -13852 4488 -13366
rect 4170 -14012 4296 -14002
rect 4802 -13134 4928 -13124
rect 4614 -13852 4802 -13366
rect 4488 -14012 4614 -14002
rect 5118 -13134 5244 -13124
rect 4928 -13852 5118 -13366
rect 4802 -14014 4928 -14004
rect 5436 -13134 5562 -13124
rect 5244 -13852 5436 -13366
rect 5118 -14014 5244 -14004
rect 5750 -13134 5876 -13124
rect 5562 -13852 5750 -13366
rect 5436 -14014 5562 -14004
rect 5750 -14014 5876 -14004
rect -4594 -14118 -4534 -14108
rect -4274 -14116 -4214 -14106
rect -4534 -14228 -4274 -14134
rect -4594 -14258 -4534 -14248
rect -4646 -14540 -4538 -14530
rect -5606 -14641 -4646 -14563
rect -4646 -14672 -4538 -14662
rect -5896 -14916 -5756 -14906
rect -4479 -14979 -4393 -14228
rect -4274 -14256 -4214 -14246
rect -3544 -14374 -3418 -14364
rect -5756 -15065 -4393 -14979
rect -4277 -15007 -4271 -14933
rect -4197 -15007 -4027 -14933
rect -5896 -15130 -5756 -15120
rect -4479 -15484 -4393 -15065
rect -4694 -15494 -4634 -15484
rect -4479 -15494 -4316 -15484
rect -4479 -15514 -4376 -15494
rect -4634 -15600 -4376 -15514
rect -4694 -15634 -4634 -15624
rect -4376 -15634 -4316 -15624
rect -5400 -16184 -5330 -16174
rect -5725 -16296 -5400 -16210
rect -5725 -18644 -5639 -16296
rect -4850 -16186 -4790 -16176
rect -5330 -16296 -4850 -16210
rect -5400 -16328 -5330 -16318
rect -4530 -16184 -4470 -16174
rect -4790 -16296 -4530 -16210
rect -4850 -16326 -4790 -16316
rect -4220 -16190 -4160 -16180
rect -4470 -16296 -4220 -16210
rect -4530 -16324 -4470 -16314
rect -4101 -16215 -4027 -15007
rect -3226 -14374 -3100 -14364
rect -3418 -15068 -3226 -14534
rect -3544 -15254 -3418 -15244
rect -2912 -14376 -2786 -14366
rect -3100 -15068 -2912 -14534
rect -3226 -15254 -3100 -15244
rect -2596 -14376 -2470 -14366
rect -2786 -15068 -2596 -14534
rect -2912 -15256 -2786 -15246
rect -2278 -14376 -2152 -14366
rect -2470 -15068 -2278 -14534
rect -2596 -15256 -2470 -15246
rect -1558 -14374 -1432 -14364
rect -2152 -15068 -1558 -14534
rect -2278 -15256 -2152 -15246
rect -1240 -14374 -1114 -14364
rect -1432 -15068 -1240 -14534
rect -1558 -15254 -1432 -15244
rect -926 -14376 -800 -14366
rect -1114 -15068 -926 -14534
rect -1240 -15254 -1114 -15244
rect -610 -14376 -484 -14366
rect -800 -15068 -610 -14534
rect -926 -15256 -800 -15246
rect -292 -14376 -166 -14366
rect -484 -15068 -292 -14534
rect -610 -15256 -484 -15246
rect 404 -14374 530 -14364
rect -166 -15068 404 -14534
rect -292 -15256 -166 -15246
rect 722 -14374 848 -14364
rect 530 -15068 722 -14534
rect 404 -15254 530 -15244
rect 1036 -14376 1162 -14366
rect 848 -15068 1036 -14534
rect 722 -15254 848 -15244
rect 1352 -14376 1478 -14366
rect 1162 -15068 1352 -14534
rect 1036 -15256 1162 -15246
rect 1670 -14376 1796 -14366
rect 1478 -15068 1670 -14534
rect 1352 -15256 1478 -15246
rect 2366 -14380 2492 -14370
rect 1796 -15068 2366 -14534
rect 1670 -15256 1796 -15246
rect 2684 -14380 2810 -14370
rect 2492 -15068 2684 -14534
rect 2366 -15260 2492 -15250
rect 2998 -14382 3124 -14372
rect 2810 -15068 2998 -14534
rect 2684 -15260 2810 -15250
rect 3314 -14382 3440 -14372
rect 3124 -15068 3314 -14534
rect 2998 -15262 3124 -15252
rect 3632 -14382 3758 -14372
rect 3440 -15068 3632 -14534
rect 3314 -15262 3440 -15252
rect 4324 -14380 4450 -14370
rect 3758 -14550 4324 -14534
rect 4642 -14380 4768 -14370
rect 4450 -14550 4642 -14534
rect 4956 -14382 5082 -14372
rect 4768 -14550 4956 -14534
rect 5272 -14382 5398 -14372
rect 5082 -14550 5272 -14534
rect 5590 -14382 5716 -14372
rect 5398 -14550 5590 -14534
rect 3758 -15060 3814 -14550
rect 3758 -15068 4324 -15060
rect 3814 -15070 4324 -15068
rect 3632 -15262 3758 -15252
rect 4450 -15070 4642 -15060
rect 4324 -15260 4450 -15250
rect 4768 -15070 4956 -15060
rect 4642 -15260 4768 -15250
rect 5082 -15070 5272 -15060
rect 4956 -15262 5082 -15252
rect 5398 -15070 5590 -15060
rect 5272 -15262 5398 -15252
rect 5590 -15262 5716 -15252
rect -4160 -16289 -4027 -16215
rect -3698 -15362 -3572 -15352
rect -3380 -15362 -3254 -15352
rect -3572 -16042 -3380 -15556
rect -3698 -16242 -3572 -16232
rect -3066 -15364 -2940 -15354
rect -3254 -15610 -3066 -15556
rect -2750 -15364 -2624 -15354
rect -2940 -15610 -2750 -15556
rect -2432 -15364 -2306 -15354
rect -2624 -15610 -2432 -15556
rect -2118 -15364 -1992 -15354
rect -2306 -15610 -2118 -15556
rect -1712 -15362 -1586 -15352
rect -1924 -15552 -1786 -15542
rect -1992 -15610 -1924 -15556
rect -1786 -15610 -1712 -15556
rect -1394 -15362 -1268 -15352
rect -1586 -15610 -1394 -15556
rect -1080 -15364 -954 -15354
rect -1268 -15610 -1080 -15556
rect -764 -15364 -638 -15354
rect -954 -15610 -764 -15556
rect -446 -15364 -320 -15354
rect -638 -15610 -446 -15556
rect -132 -15364 -6 -15354
rect -320 -15610 -132 -15556
rect -3254 -15924 -3202 -15610
rect -3254 -16042 -3066 -15924
rect -3380 -16242 -3254 -16232
rect -2940 -16042 -2750 -15924
rect -3066 -16244 -2940 -16234
rect -2624 -16042 -2432 -15924
rect -2750 -16244 -2624 -16234
rect -2306 -16042 -2118 -15924
rect -2432 -16244 -2306 -16234
rect -1992 -16036 -1924 -15924
rect -1786 -16036 -1712 -15924
rect -1992 -16042 -1712 -16036
rect -1924 -16046 -1786 -16042
rect -2118 -16244 -1992 -16234
rect -1586 -16042 -1394 -15924
rect -1712 -16242 -1586 -16232
rect -1268 -16042 -1080 -15924
rect -1394 -16242 -1268 -16232
rect -954 -16042 -764 -15924
rect -1080 -16244 -954 -16234
rect -638 -16042 -446 -15924
rect -764 -16244 -638 -16234
rect -320 -16042 -132 -15924
rect -446 -16244 -320 -16234
rect 250 -15362 376 -15352
rect -6 -15610 250 -15556
rect -6 -16042 250 -15924
rect -132 -16244 -6 -16234
rect 568 -15362 694 -15352
rect 376 -15610 568 -15556
rect 376 -16042 568 -15924
rect 250 -16242 376 -16232
rect 882 -15364 1008 -15354
rect 694 -15610 882 -15556
rect 694 -16042 882 -15924
rect 568 -16242 694 -16232
rect 1198 -15364 1324 -15354
rect 1008 -15610 1198 -15556
rect 1008 -16042 1198 -15924
rect 882 -16244 1008 -16234
rect 1516 -15364 1642 -15354
rect 1324 -15610 1516 -15556
rect 1324 -16042 1516 -15924
rect 1198 -16244 1324 -16234
rect 1830 -15364 1956 -15354
rect 1642 -15610 1830 -15556
rect 1642 -16042 1830 -15924
rect 1516 -16244 1642 -16234
rect 2212 -15368 2338 -15358
rect 2022 -15556 2160 -15550
rect 1956 -15560 2212 -15556
rect 1956 -15610 2022 -15560
rect 1956 -16042 2022 -15924
rect 2160 -15610 2212 -15560
rect 2160 -16042 2212 -15924
rect 2022 -16054 2160 -16044
rect 1830 -16244 1956 -16234
rect 2530 -15368 2656 -15358
rect 2338 -15610 2530 -15556
rect 2338 -16042 2530 -15924
rect 2212 -16248 2338 -16238
rect 2844 -15370 2970 -15360
rect 2656 -15610 2844 -15556
rect 2656 -16042 2844 -15924
rect 2530 -16248 2656 -16238
rect 3160 -15370 3286 -15360
rect 2970 -15610 3160 -15556
rect 2970 -16042 3160 -15924
rect 2844 -16250 2970 -16240
rect 3478 -15370 3604 -15360
rect 3286 -15610 3478 -15556
rect 3332 -15924 3478 -15610
rect 3286 -16042 3478 -15924
rect 3160 -16250 3286 -16240
rect 3792 -15370 3918 -15360
rect 3604 -16042 3792 -15556
rect 3478 -16250 3604 -16240
rect 4170 -15368 4296 -15358
rect 3918 -16042 4170 -15556
rect 3792 -16250 3918 -16240
rect 4488 -15368 4614 -15358
rect 4296 -16042 4488 -15556
rect 4170 -16248 4296 -16238
rect 4802 -15370 4928 -15360
rect 4614 -16042 4802 -15556
rect 4488 -16248 4614 -16238
rect 5118 -15370 5244 -15360
rect 4928 -16042 5118 -15556
rect 4802 -16250 4928 -16240
rect 5436 -15370 5562 -15360
rect 5244 -16042 5436 -15556
rect 5118 -16250 5244 -16240
rect 5750 -15370 5876 -15360
rect 5562 -16042 5750 -15556
rect 5436 -16250 5562 -16240
rect 5750 -16250 5876 -16240
rect -4220 -16330 -4160 -16320
rect -3908 -16912 -3786 -16902
rect -5542 -16994 -5482 -16984
rect -5228 -16994 -5168 -16984
rect -5482 -17112 -5228 -17006
rect -5542 -17134 -5482 -17124
rect -4912 -16996 -4852 -16986
rect -5168 -17112 -4912 -17006
rect -5228 -17134 -5168 -17124
rect -4594 -16996 -4534 -16986
rect -4852 -17112 -4594 -17006
rect -4912 -17136 -4852 -17126
rect -4276 -16998 -4216 -16988
rect -4534 -17112 -4276 -17006
rect -4594 -17136 -4534 -17126
rect -4216 -17112 -3908 -17006
rect -4276 -17138 -4216 -17128
rect -3908 -17180 -3786 -17170
rect -3544 -16980 -3418 -16970
rect -3226 -16980 -3100 -16970
rect -3418 -17668 -3226 -17134
rect -3544 -17860 -3418 -17850
rect -2912 -16982 -2786 -16972
rect -3100 -17668 -2912 -17134
rect -3226 -17860 -3100 -17850
rect -2596 -16982 -2470 -16972
rect -2786 -17668 -2596 -17134
rect -2912 -17862 -2786 -17852
rect -2278 -16982 -2152 -16972
rect -2470 -17668 -2278 -17134
rect -2596 -17862 -2470 -17852
rect -1558 -16980 -1432 -16970
rect -2152 -17668 -1558 -17134
rect -2278 -17862 -2152 -17852
rect -1240 -16980 -1114 -16970
rect -1432 -17668 -1240 -17134
rect -1558 -17860 -1432 -17850
rect -926 -16982 -800 -16972
rect -1114 -17668 -926 -17134
rect -1240 -17860 -1114 -17850
rect -610 -16982 -484 -16972
rect -800 -17668 -610 -17134
rect -926 -17862 -800 -17852
rect -292 -16982 -166 -16972
rect -484 -17668 -292 -17134
rect -610 -17862 -484 -17852
rect 404 -16980 530 -16970
rect -166 -17668 404 -17134
rect -292 -17862 -166 -17852
rect 722 -16980 848 -16970
rect 530 -17668 722 -17134
rect 404 -17860 530 -17850
rect 1036 -16982 1162 -16972
rect 848 -17668 1036 -17134
rect 722 -17860 848 -17850
rect 1352 -16982 1478 -16972
rect 1162 -17668 1352 -17134
rect 1036 -17862 1162 -17852
rect 1670 -16982 1796 -16972
rect 1478 -17668 1670 -17134
rect 1352 -17862 1478 -17852
rect 2366 -16986 2492 -16976
rect 1796 -17668 2366 -17134
rect 1670 -17862 1796 -17852
rect 2684 -16986 2810 -16976
rect 2492 -17668 2684 -17134
rect 2366 -17866 2492 -17856
rect 2998 -16988 3124 -16978
rect 2810 -17668 2998 -17134
rect 2684 -17866 2810 -17856
rect 3314 -16988 3440 -16978
rect 3124 -17668 3314 -17134
rect 2998 -17868 3124 -17858
rect 3632 -16988 3758 -16978
rect 3440 -17668 3632 -17134
rect 3314 -17868 3440 -17858
rect 4324 -16986 4450 -16976
rect 3810 -17134 4324 -17130
rect 3758 -17140 4324 -17134
rect 4642 -16986 4768 -16976
rect 4450 -17140 4642 -17130
rect 4956 -16988 5082 -16978
rect 4768 -17140 4956 -17130
rect 5272 -16988 5398 -16978
rect 5082 -17140 5272 -17130
rect 5590 -16988 5716 -16978
rect 5398 -17140 5590 -17130
rect 3758 -17650 3810 -17140
rect 3758 -17668 4324 -17650
rect 3632 -17868 3758 -17858
rect 4450 -17668 4642 -17650
rect 4324 -17866 4450 -17856
rect 4768 -17668 4956 -17650
rect 4642 -17866 4768 -17856
rect 5082 -17668 5272 -17650
rect 4956 -17868 5082 -17858
rect 5398 -17668 5590 -17650
rect 5272 -17868 5398 -17858
rect 5590 -17868 5716 -17858
rect -3698 -17968 -3572 -17958
rect -5725 -18774 -5702 -18644
rect -5642 -18670 -5639 -18644
rect -5386 -18646 -5326 -18636
rect -5642 -18762 -5386 -18670
rect -5642 -18774 -5639 -18762
rect -5725 -18791 -5639 -18774
rect -5068 -18646 -5008 -18636
rect -5326 -18762 -5068 -18670
rect -5386 -18786 -5326 -18776
rect -4752 -18646 -4692 -18636
rect -5008 -18762 -4752 -18670
rect -5068 -18786 -5008 -18776
rect -4436 -18646 -4376 -18636
rect -4692 -18762 -4436 -18670
rect -4752 -18786 -4692 -18776
rect -4118 -18646 -4058 -18636
rect -4376 -18762 -4118 -18670
rect -4436 -18786 -4376 -18776
rect -4058 -18762 -3698 -18670
rect -4118 -18786 -4058 -18776
rect -3380 -17968 -3254 -17958
rect -3572 -18652 -3380 -18166
rect -3698 -18848 -3572 -18838
rect -3066 -17970 -2940 -17960
rect -3254 -18652 -3066 -18166
rect -3380 -18848 -3254 -18838
rect -2750 -17970 -2624 -17960
rect -2940 -18652 -2750 -18166
rect -3066 -18850 -2940 -18840
rect -2432 -17970 -2306 -17960
rect -2624 -18652 -2432 -18166
rect -2750 -18850 -2624 -18840
rect -2118 -17970 -1992 -17960
rect -2306 -18652 -2118 -18166
rect -2432 -18850 -2306 -18840
rect -1712 -17968 -1586 -17958
rect -1992 -18652 -1712 -18166
rect -2118 -18850 -1992 -18840
rect -1394 -17968 -1268 -17958
rect -1586 -18652 -1394 -18166
rect -1712 -18848 -1586 -18838
rect -1080 -17970 -954 -17960
rect -1268 -18652 -1080 -18166
rect -1394 -18848 -1268 -18838
rect -764 -17970 -638 -17960
rect -954 -18652 -764 -18166
rect -1080 -18850 -954 -18840
rect -446 -17970 -320 -17960
rect -638 -18652 -446 -18166
rect -764 -18850 -638 -18840
rect -132 -17970 -6 -17960
rect -320 -18652 -132 -18166
rect -446 -18850 -320 -18840
rect 250 -17968 376 -17958
rect 56 -18164 194 -18154
rect -6 -18320 56 -18166
rect 194 -18320 250 -18166
rect 568 -17968 694 -17958
rect 376 -18320 568 -18166
rect 882 -17970 1008 -17960
rect 694 -18320 882 -18166
rect 1198 -17970 1324 -17960
rect 1008 -18320 1198 -18166
rect 1516 -17970 1642 -17960
rect 1324 -18320 1516 -18166
rect 1830 -17970 1956 -17960
rect 1642 -18320 1830 -18166
rect 2212 -17974 2338 -17964
rect 1956 -18320 2212 -18166
rect 2530 -17974 2656 -17964
rect 2338 -18320 2530 -18166
rect 2844 -17976 2970 -17966
rect 2656 -18320 2844 -18166
rect 3160 -17976 3286 -17966
rect 2970 -18320 3160 -18166
rect 3478 -17976 3604 -17966
rect -6 -18634 34 -18320
rect -6 -18648 56 -18634
rect 194 -18648 250 -18634
rect -6 -18652 250 -18648
rect 56 -18658 194 -18652
rect -132 -18850 -6 -18840
rect 376 -18652 568 -18634
rect 250 -18848 376 -18838
rect 694 -18652 882 -18634
rect 568 -18848 694 -18838
rect 1008 -18652 1198 -18634
rect 882 -18850 1008 -18840
rect 1324 -18652 1516 -18634
rect 1198 -18850 1324 -18840
rect 1642 -18652 1830 -18634
rect 1516 -18850 1642 -18840
rect 1956 -18652 2212 -18634
rect 1830 -18850 1956 -18840
rect 2338 -18652 2530 -18634
rect 2212 -18854 2338 -18844
rect 2656 -18652 2844 -18634
rect 2530 -18854 2656 -18844
rect 2970 -18652 3160 -18634
rect 2844 -18856 2970 -18846
rect 3286 -18652 3478 -18166
rect 3160 -18856 3286 -18846
rect 3792 -17976 3918 -17966
rect 3604 -18652 3792 -18166
rect 3478 -18856 3604 -18846
rect 4170 -17974 4296 -17964
rect 3972 -18164 4110 -18154
rect 3918 -18648 3972 -18166
rect 4110 -18648 4170 -18166
rect 3918 -18652 4170 -18648
rect 3972 -18658 4110 -18652
rect 3792 -18856 3918 -18846
rect 4488 -17974 4614 -17964
rect 4296 -18652 4488 -18166
rect 4170 -18854 4296 -18844
rect 4802 -17976 4928 -17966
rect 4614 -18652 4802 -18166
rect 4488 -18854 4614 -18844
rect 5118 -17976 5244 -17966
rect 4928 -18652 5118 -18166
rect 4802 -18856 4928 -18846
rect 5436 -17976 5562 -17966
rect 5244 -18652 5436 -18166
rect 5118 -18856 5244 -18846
rect 5750 -17976 5876 -17966
rect 5562 -18652 5750 -18166
rect 5436 -18856 5562 -18846
rect 5750 -18856 5876 -18846
rect -3542 -19190 -3416 -19180
rect -3224 -19190 -3098 -19180
rect -3416 -19918 -3224 -19384
rect -3542 -20070 -3416 -20060
rect -2910 -19192 -2784 -19182
rect -3098 -19918 -2910 -19384
rect -3224 -20070 -3098 -20060
rect -2594 -19192 -2468 -19182
rect -2784 -19918 -2594 -19384
rect -2910 -20072 -2784 -20062
rect -2276 -19192 -2150 -19182
rect -2468 -19918 -2276 -19384
rect -2594 -20072 -2468 -20062
rect -1556 -19190 -1430 -19180
rect -2150 -19918 -1556 -19384
rect -2276 -20072 -2150 -20062
rect -1238 -19190 -1112 -19180
rect -1430 -19918 -1238 -19384
rect -1556 -20070 -1430 -20060
rect -924 -19192 -798 -19182
rect -1112 -19918 -924 -19384
rect -1238 -20070 -1112 -20060
rect -608 -19192 -482 -19182
rect -798 -19918 -608 -19384
rect -924 -20072 -798 -20062
rect -290 -19192 -164 -19182
rect -482 -19918 -290 -19384
rect -608 -20072 -482 -20062
rect 406 -19190 532 -19180
rect -164 -19918 406 -19384
rect -290 -20072 -164 -20062
rect 724 -19190 850 -19180
rect 532 -19918 724 -19384
rect 406 -20070 532 -20060
rect 1038 -19192 1164 -19182
rect 850 -19918 1038 -19384
rect 724 -20070 850 -20060
rect 1354 -19192 1480 -19182
rect 1164 -19918 1354 -19384
rect 1038 -20072 1164 -20062
rect 1672 -19192 1798 -19182
rect 1480 -19918 1672 -19384
rect 1354 -20072 1480 -20062
rect 2368 -19196 2494 -19186
rect 1798 -19918 2368 -19384
rect 1672 -20072 1798 -20062
rect 2686 -19196 2812 -19186
rect 2494 -19918 2686 -19384
rect 2368 -20076 2494 -20066
rect 3000 -19198 3126 -19188
rect 2812 -19918 3000 -19384
rect 2686 -20076 2812 -20066
rect 3316 -19198 3442 -19188
rect 3126 -19918 3316 -19384
rect 3000 -20078 3126 -20068
rect 3634 -19198 3760 -19188
rect 3442 -19918 3634 -19384
rect 3316 -20078 3442 -20068
rect 4326 -19196 4452 -19186
rect 3760 -19400 4326 -19384
rect 4644 -19196 4770 -19186
rect 4452 -19400 4644 -19384
rect 4958 -19198 5084 -19188
rect 4770 -19400 4958 -19384
rect 5274 -19198 5400 -19188
rect 5084 -19400 5274 -19384
rect 5592 -19198 5718 -19188
rect 5400 -19400 5592 -19384
rect 3760 -19910 3808 -19400
rect 3760 -19918 4326 -19910
rect 3808 -19920 4326 -19918
rect 3634 -20078 3760 -20068
rect 4452 -19920 4644 -19910
rect 4326 -20076 4452 -20066
rect 4770 -19920 4958 -19910
rect 4644 -20076 4770 -20066
rect 5084 -19920 5274 -19910
rect 4958 -20078 5084 -20068
rect 5400 -19920 5592 -19910
rect 5274 -20078 5400 -20068
rect 5592 -20078 5718 -20068
rect -3696 -20178 -3570 -20168
rect -3378 -20178 -3252 -20168
rect -3570 -20874 -3378 -20388
rect -3696 -21058 -3570 -21048
rect -3064 -20180 -2938 -20170
rect -3252 -20874 -3064 -20388
rect -3378 -21058 -3252 -21048
rect -2748 -20180 -2622 -20170
rect -2938 -20874 -2748 -20388
rect -3064 -21060 -2938 -21050
rect -2430 -20180 -2304 -20170
rect -2622 -20874 -2430 -20388
rect -2748 -21060 -2622 -21050
rect -2116 -20180 -1990 -20170
rect -2304 -20874 -2116 -20388
rect -2430 -21060 -2304 -21050
rect -1710 -20178 -1584 -20168
rect -1918 -20388 -1780 -20380
rect -1990 -20390 -1710 -20388
rect -1990 -20874 -1918 -20390
rect -1780 -20874 -1710 -20390
rect -1918 -20884 -1780 -20874
rect -2116 -21060 -1990 -21050
rect -1392 -20178 -1266 -20168
rect -1584 -20874 -1392 -20388
rect -1710 -21058 -1584 -21048
rect -1078 -20180 -952 -20170
rect -1266 -20874 -1078 -20388
rect -1392 -21058 -1266 -21048
rect -762 -20180 -636 -20170
rect -952 -20874 -762 -20388
rect -1078 -21060 -952 -21050
rect -444 -20180 -318 -20170
rect -636 -20874 -444 -20388
rect -762 -21060 -636 -21050
rect -130 -20180 -4 -20170
rect -318 -20874 -130 -20388
rect -444 -21060 -318 -21050
rect 252 -20178 378 -20168
rect -4 -20468 252 -20388
rect 570 -20178 696 -20168
rect 378 -20468 570 -20388
rect 884 -20180 1010 -20170
rect 696 -20468 884 -20388
rect 1200 -20180 1326 -20170
rect 1010 -20468 1200 -20388
rect 1518 -20180 1644 -20170
rect 1326 -20468 1518 -20388
rect 1832 -20180 1958 -20170
rect 1644 -20468 1832 -20388
rect 2214 -20184 2340 -20174
rect 2016 -20388 2154 -20378
rect 1958 -20468 2016 -20388
rect 2154 -20468 2214 -20388
rect 2532 -20184 2658 -20174
rect 2340 -20468 2532 -20388
rect 2846 -20186 2972 -20176
rect 2658 -20468 2846 -20388
rect 3162 -20186 3288 -20176
rect 2972 -20468 3162 -20388
rect 3480 -20186 3606 -20176
rect -4 -20782 52 -20468
rect -4 -20874 252 -20782
rect -130 -21060 -4 -21050
rect 378 -20874 570 -20782
rect 252 -21058 378 -21048
rect 696 -20874 884 -20782
rect 570 -21058 696 -21048
rect 1010 -20874 1200 -20782
rect 884 -21060 1010 -21050
rect 1326 -20874 1518 -20782
rect 1200 -21060 1326 -21050
rect 1644 -20874 1832 -20782
rect 1518 -21060 1644 -21050
rect 1958 -20872 2016 -20782
rect 2154 -20872 2214 -20782
rect 1958 -20874 2214 -20872
rect 2016 -20882 2154 -20874
rect 1832 -21060 1958 -21050
rect 2340 -20874 2532 -20782
rect 2214 -21064 2340 -21054
rect 2658 -20874 2846 -20782
rect 2532 -21064 2658 -21054
rect 2972 -20874 3162 -20782
rect 2846 -21066 2972 -21056
rect 3288 -20874 3480 -20388
rect 3162 -21066 3288 -21056
rect 3794 -20186 3920 -20176
rect 3606 -20874 3794 -20388
rect 3480 -21066 3606 -21056
rect 4172 -20184 4298 -20174
rect 3920 -20874 4172 -20388
rect 3794 -21066 3920 -21056
rect 4490 -20184 4616 -20174
rect 4298 -20874 4490 -20388
rect 4172 -21064 4298 -21054
rect 4804 -20186 4930 -20176
rect 4616 -20874 4804 -20388
rect 4490 -21064 4616 -21054
rect 5120 -20186 5246 -20176
rect 4930 -20874 5120 -20388
rect 4804 -21066 4930 -21056
rect 5438 -20186 5564 -20176
rect 5246 -20874 5438 -20388
rect 5120 -21066 5246 -21056
rect 5752 -20186 5878 -20176
rect 5564 -20874 5752 -20388
rect 5438 -21066 5564 -21056
rect 5752 -21066 5878 -21056
<< via2 >>
rect 3808 -8356 4324 -7846
rect 4324 -8356 4450 -7846
rect 4450 -8356 4642 -7846
rect 4642 -8356 4768 -7846
rect 4768 -8356 4956 -7846
rect 4956 -8356 5082 -7846
rect 5082 -8356 5272 -7846
rect 5272 -8356 5398 -7846
rect 5398 -8356 5590 -7846
rect 5590 -8356 5628 -7846
rect -3202 -9336 -3066 -9022
rect -3066 -9336 -2940 -9022
rect -2940 -9336 -2750 -9022
rect -2750 -9336 -2624 -9022
rect -2624 -9336 -2432 -9022
rect -2432 -9336 -2306 -9022
rect -2306 -9336 -2118 -9022
rect -2118 -9336 -1992 -9022
rect -1992 -9336 -1712 -9022
rect -1712 -9336 -1586 -9022
rect -1586 -9336 -1394 -9022
rect -1394 -9336 -1268 -9022
rect -1268 -9336 -1080 -9022
rect -1080 -9336 -954 -9022
rect -954 -9336 -764 -9022
rect -764 -9336 -638 -9022
rect -638 -9336 -446 -9022
rect -446 -9336 -320 -9022
rect -320 -9336 -208 -9022
rect 3808 -10602 4324 -10092
rect 4324 -10602 4450 -10092
rect 4450 -10602 4642 -10092
rect 4642 -10602 4768 -10092
rect 4768 -10602 4956 -10092
rect 4956 -10602 5082 -10092
rect 5082 -10602 5272 -10092
rect 5272 -10602 5398 -10092
rect 5398 -10602 5590 -10092
rect 5590 -10602 5628 -10092
rect -3214 -11548 -3066 -11234
rect -3066 -11548 -2940 -11234
rect -2940 -11548 -2750 -11234
rect -2750 -11548 -2624 -11234
rect -2624 -11548 -2432 -11234
rect -2432 -11548 -2306 -11234
rect -2306 -11548 -2118 -11234
rect -2118 -11548 -1992 -11234
rect -1992 -11548 -1920 -11234
rect -1920 -11548 -1782 -11234
rect -1782 -11548 -1712 -11234
rect -1712 -11548 -1586 -11234
rect -1586 -11548 -1394 -11234
rect -1394 -11548 -1268 -11234
rect -1268 -11548 -1080 -11234
rect -1080 -11548 -954 -11234
rect -954 -11548 -764 -11234
rect -764 -11548 -638 -11234
rect -638 -11548 -446 -11234
rect -446 -11548 -320 -11234
rect -320 -11548 -176 -11234
rect 3808 -12794 4324 -12284
rect 4324 -12794 4450 -12284
rect 4450 -12794 4642 -12284
rect 4642 -12794 4768 -12284
rect 4768 -12794 4956 -12284
rect 4956 -12794 5082 -12284
rect 5082 -12794 5272 -12284
rect 5272 -12794 5398 -12284
rect 5398 -12794 5590 -12284
rect 5590 -12794 5628 -12284
rect -3208 -13802 -3066 -13488
rect -3066 -13802 -2940 -13488
rect -2940 -13802 -2750 -13488
rect -2750 -13802 -2624 -13488
rect -2624 -13802 -2432 -13488
rect -2432 -13802 -2306 -13488
rect -2306 -13802 -2118 -13488
rect -2118 -13802 -1992 -13488
rect -1992 -13802 -1712 -13488
rect -1712 -13802 -1586 -13488
rect -1586 -13802 -1394 -13488
rect -1394 -13802 -1268 -13488
rect -1268 -13802 -1080 -13488
rect -1080 -13802 -954 -13488
rect -954 -13802 -764 -13488
rect -764 -13802 -638 -13488
rect -638 -13802 -446 -13488
rect -446 -13802 -320 -13488
rect -320 -13802 -194 -13488
rect 3814 -15060 4324 -14550
rect 4324 -15060 4450 -14550
rect 4450 -15060 4642 -14550
rect 4642 -15060 4768 -14550
rect 4768 -15060 4956 -14550
rect 4956 -15060 5082 -14550
rect 5082 -15060 5272 -14550
rect 5272 -15060 5398 -14550
rect 5398 -15060 5590 -14550
rect 5590 -15060 5634 -14550
rect -3202 -15924 -3066 -15610
rect -3066 -15924 -2940 -15610
rect -2940 -15924 -2750 -15610
rect -2750 -15924 -2624 -15610
rect -2624 -15924 -2432 -15610
rect -2432 -15924 -2306 -15610
rect -2306 -15924 -2118 -15610
rect -2118 -15924 -1992 -15610
rect -1992 -15924 -1924 -15610
rect -1924 -15924 -1786 -15610
rect -1786 -15924 -1712 -15610
rect -1712 -15924 -1586 -15610
rect -1586 -15924 -1394 -15610
rect -1394 -15924 -1268 -15610
rect -1268 -15924 -1080 -15610
rect -1080 -15924 -954 -15610
rect -954 -15924 -764 -15610
rect -764 -15924 -638 -15610
rect -638 -15924 -446 -15610
rect -446 -15924 -320 -15610
rect -320 -15924 -165 -15610
rect 3810 -17650 4324 -17140
rect 4324 -17650 4450 -17140
rect 4450 -17650 4642 -17140
rect 4642 -17650 4768 -17140
rect 4768 -17650 4956 -17140
rect 4956 -17650 5082 -17140
rect 5082 -17650 5272 -17140
rect 5272 -17650 5398 -17140
rect 5398 -17650 5590 -17140
rect 5590 -17650 5630 -17140
rect 34 -18634 56 -18320
rect 56 -18634 194 -18320
rect 194 -18634 250 -18320
rect 250 -18634 376 -18320
rect 376 -18634 568 -18320
rect 568 -18634 694 -18320
rect 694 -18634 882 -18320
rect 882 -18634 1008 -18320
rect 1008 -18634 1198 -18320
rect 1198 -18634 1324 -18320
rect 1324 -18634 1516 -18320
rect 1516 -18634 1642 -18320
rect 1642 -18634 1830 -18320
rect 1830 -18634 1956 -18320
rect 1956 -18634 2212 -18320
rect 2212 -18634 2338 -18320
rect 2338 -18634 2530 -18320
rect 2530 -18634 2656 -18320
rect 2656 -18634 2844 -18320
rect 2844 -18634 2970 -18320
rect 2970 -18634 3160 -18320
rect 3160 -18634 3266 -18320
rect 3808 -19910 4326 -19400
rect 4326 -19910 4452 -19400
rect 4452 -19910 4644 -19400
rect 4644 -19910 4770 -19400
rect 4770 -19910 4958 -19400
rect 4958 -19910 5084 -19400
rect 5084 -19910 5274 -19400
rect 5274 -19910 5400 -19400
rect 5400 -19910 5592 -19400
rect 5592 -19910 5628 -19400
rect 52 -20782 252 -20468
rect 252 -20782 378 -20468
rect 378 -20782 570 -20468
rect 570 -20782 696 -20468
rect 696 -20782 884 -20468
rect 884 -20782 1010 -20468
rect 1010 -20782 1200 -20468
rect 1200 -20782 1326 -20468
rect 1326 -20782 1518 -20468
rect 1518 -20782 1644 -20468
rect 1644 -20782 1832 -20468
rect 1832 -20782 1958 -20468
rect 1958 -20782 2016 -20468
rect 2016 -20782 2154 -20468
rect 2154 -20782 2214 -20468
rect 2214 -20782 2340 -20468
rect 2340 -20782 2532 -20468
rect 2532 -20782 2658 -20468
rect 2658 -20782 2846 -20468
rect 2846 -20782 2972 -20468
rect 2972 -20782 3162 -20468
rect 3162 -20782 3278 -20468
<< metal3 >>
rect 3798 -7846 5638 -7841
rect 3798 -8356 3808 -7846
rect 5628 -7876 5638 -7846
rect 5628 -8356 5640 -7876
rect 3798 -8361 5640 -8356
rect -3244 -9022 -160 -8966
rect -3244 -9336 -3202 -9022
rect -208 -9336 -160 -9022
rect -3244 -11234 -160 -9336
rect 3804 -10087 5640 -8361
rect 3798 -10092 5640 -10087
rect 3798 -10602 3808 -10092
rect 5628 -10602 5640 -10092
rect 3798 -10607 5640 -10602
rect -3244 -11548 -3214 -11234
rect -176 -11548 -160 -11234
rect -3244 -13488 -160 -11548
rect 3804 -12279 5640 -10607
rect 3798 -12284 5640 -12279
rect 3798 -12794 3808 -12284
rect 5628 -12794 5640 -12284
rect 3798 -12799 5640 -12794
rect -3244 -13802 -3208 -13488
rect -194 -13802 -160 -13488
rect -3244 -15610 -160 -13802
rect -3244 -15924 -3202 -15610
rect -165 -15924 -160 -15610
rect -3244 -15966 -160 -15924
rect 3804 -14545 5640 -12799
rect 3804 -14550 5644 -14545
rect 3804 -15060 3814 -14550
rect 5634 -15060 5644 -14550
rect 3804 -15065 5644 -15060
rect 3804 -17135 5640 -15065
rect 3800 -17140 5640 -17135
rect 3800 -17650 3810 -17140
rect 5630 -17650 5640 -17140
rect 3800 -17655 5640 -17650
rect 26 -18320 3354 -18310
rect 26 -18634 34 -18320
rect 3266 -18634 3354 -18320
rect 26 -20468 3354 -18634
rect 3804 -19395 5640 -17655
rect 3798 -19400 5640 -19395
rect 3798 -19910 3808 -19400
rect 5628 -19886 5640 -19400
rect 5628 -19910 5638 -19886
rect 3798 -19915 5638 -19910
rect 26 -20782 52 -20468
rect 3278 -20782 3354 -20468
rect 26 -20810 3354 -20782
use sky130_fd_pr__nfet_g5v0d10v5_8WF6SK  sky130_fd_pr__nfet_g5v0d10v5_8WF6SK_1
timestamp 1644523392
transform 1 0 -4881 0 1 -17890
box -988 -1258 988 1258
use sky130_fd_pr__nfet_g5v0d10v5_GYVFE6  sky130_fd_pr__nfet_g5v0d10v5_GYVFE6_0
timestamp 1644523392
transform 1 0 1105 0 1 -18995
box -988 -2366 988 2366
use sky130_fd_pr__nfet_g5v0d10v5_GYVFE6  sky130_fd_pr__nfet_g5v0d10v5_GYVFE6_1
timestamp 1644523392
transform 1 0 -855 0 1 -18995
box -988 -2366 988 2366
use sky130_fd_pr__nfet_g5v0d10v5_GYVFE6  sky130_fd_pr__nfet_g5v0d10v5_GYVFE6_2
timestamp 1644523392
transform 1 0 -2843 0 1 -18995
box -988 -2366 988 2366
use sky130_fd_pr__nfet_g5v0d10v5_GYVFE6  sky130_fd_pr__nfet_g5v0d10v5_GYVFE6_3
timestamp 1644523392
transform 1 0 5025 0 1 -18995
box -988 -2366 988 2366
use sky130_fd_pr__nfet_g5v0d10v5_GYVFE6  sky130_fd_pr__nfet_g5v0d10v5_GYVFE6_4
timestamp 1644523392
transform 1 0 3065 0 1 -18995
box -988 -2366 988 2366
use sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3  sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3_0
timestamp 1644523392
transform 1 0 -5280 0 1 -15988
box -278 -658 278 658
use sky130_fd_pr__nfet_g5v0d10v5_QABAEG  sky130_fd_pr__nfet_g5v0d10v5_QABAEG_0
timestamp 1644523392
transform 1 0 -4505 0 1 -15888
box -514 -758 514 758
use sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ  sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ_0
timestamp 1644523392
transform 1 0 -5280 0 1 -14990
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_3QQKN5  sky130_fd_pr__pfet_g5v0d10v5_3QQKN5_1
timestamp 1644523392
transform 1 0 -5262 0 1 -12726
box -386 -696 386 696
use sky130_fd_pr__pfet_g5v0d10v5_CYK6CA  sky130_fd_pr__pfet_g5v0d10v5_CYK6CA_0
timestamp 1644523392
transform 1 0 1105 0 1 -11927
box -1019 -4651 1019 4651
use sky130_fd_pr__pfet_g5v0d10v5_CYK6CA  sky130_fd_pr__pfet_g5v0d10v5_CYK6CA_1
timestamp 1644523392
transform 1 0 -855 0 1 -11927
box -1019 -4651 1019 4651
use sky130_fd_pr__pfet_g5v0d10v5_CYK6CA  sky130_fd_pr__pfet_g5v0d10v5_CYK6CA_2
timestamp 1644523392
transform 1 0 -2843 0 1 -11927
box -1019 -4651 1019 4651
use sky130_fd_pr__pfet_g5v0d10v5_CYK6CA  sky130_fd_pr__pfet_g5v0d10v5_CYK6CA_3
timestamp 1644523392
transform 1 0 5025 0 1 -11927
box -1019 -4651 1019 4651
use sky130_fd_pr__pfet_g5v0d10v5_CYK6CA  sky130_fd_pr__pfet_g5v0d10v5_CYK6CA_4
timestamp 1644523392
transform 1 0 3065 0 1 -11927
box -1019 -4651 1019 4651
use sky130_fd_pr__pfet_g5v0d10v5_CYU7F7  sky130_fd_pr__pfet_g5v0d10v5_CYU7F7_0
timestamp 1644523392
transform 1 0 -4881 0 1 -9691
box -1018 -2414 1018 2414
use sky130_fd_pr__pfet_g5v0d10v5_HKUKAU  sky130_fd_pr__pfet_g5v0d10v5_HKUKAU_0
timestamp 1644523392
transform 1 0 -5263 0 1 -13774
box -386 -362 386 362
use sky130_fd_pr__pfet_g5v0d10v5_WECJAU  sky130_fd_pr__pfet_g5v0d10v5_WECJAU_0
timestamp 1644523392
transform 1 0 -4407 0 1 -13325
box -544 -1296 544 1296
<< labels >>
rlabel metal1 -5328 -14860 -5220 -13880 1 in
port 1 n
rlabel metal1 -5612 -15558 -5560 -13166 1 drv1
rlabel metal2 -5606 -14641 -4646 -14563 1 drv2
rlabel metal1 -5902 -16858 -5742 -15120 1 crosscon
port 2 n
rlabel metal1 -3923 -16912 -3769 -9948 1 drv4
rlabel metal3 3804 -14550 5640 -12794 1 out
port 3 n
rlabel metal3 26 -20468 3354 -18634 1 vss
port 5 n
rlabel metal3 -3244 -15610 -160 -13802 1 vdd_hi
port 4 n
<< end >>
