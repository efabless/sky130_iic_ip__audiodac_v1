magic
tech sky130A
magscale 1 2
timestamp 1644660372
<< mvndiff >>
rect -3307 -18881 -3273 -18869
<< locali >>
rect -814 -16844 -798 -16810
rect -3344 -19246 -930 -19060
<< viali >>
rect -2162 -15974 -2108 -15854
rect -2164 -19784 -2108 -19660
<< metal1 >>
rect -2168 -15854 -2102 -15842
rect -3098 -15974 -3088 -15854
rect -3030 -15974 -3020 -15854
rect -2782 -15974 -2772 -15854
rect -2714 -15974 -2704 -15854
rect -2466 -15974 -2456 -15854
rect -2398 -15974 -2388 -15854
rect -2172 -15974 -2162 -15854
rect -2108 -15974 -2098 -15854
rect -1882 -15974 -1872 -15854
rect -1814 -15974 -1804 -15854
rect -1566 -15974 -1556 -15854
rect -1498 -15974 -1488 -15854
rect -1250 -15974 -1240 -15854
rect -1182 -15974 -1172 -15854
rect -2168 -15986 -2102 -15974
rect -2940 -16254 -2930 -16134
rect -2872 -16254 -2862 -16134
rect -2624 -16254 -2614 -16134
rect -2556 -16254 -2546 -16134
rect -2308 -16254 -2298 -16134
rect -2240 -16254 -2230 -16134
rect -2040 -16180 -2030 -16134
rect -2146 -16254 -2030 -16180
rect -1972 -16254 -1962 -16134
rect -1724 -16254 -1714 -16134
rect -1656 -16254 -1646 -16134
rect -1408 -16254 -1398 -16134
rect -1340 -16254 -1330 -16134
rect -2146 -16256 -1962 -16254
rect -2146 -16294 -2074 -16256
rect -3026 -16342 -2074 -16294
rect -1968 -16342 -1244 -16294
rect -1968 -16372 -1896 -16342
rect -1968 -16424 -1962 -16372
rect -1910 -16424 -1896 -16372
rect -3255 -16749 -802 -16748
rect -3727 -16850 -802 -16749
rect -3727 -16851 -3255 -16850
rect -3727 -18914 -3625 -16851
rect -3570 -17222 -3560 -16990
rect -3498 -17222 -3488 -16990
rect -3092 -17222 -3082 -16990
rect -3020 -17222 -3010 -16990
rect -2616 -17222 -2606 -16990
rect -2544 -17222 -2534 -16990
rect -1760 -17222 -1750 -16990
rect -1688 -17222 -1678 -16990
rect -1284 -17222 -1274 -16990
rect -1212 -17222 -1202 -16990
rect -808 -17222 -798 -16990
rect -736 -17222 -726 -16990
rect -3326 -18882 -3316 -18804
rect -3264 -18882 -3254 -18804
rect -2850 -18882 -2840 -18804
rect -2788 -18882 -2778 -18804
rect -2374 -18882 -2364 -18804
rect -2312 -18882 -2302 -18804
rect -1994 -18882 -1984 -18804
rect -1932 -18882 -1922 -18804
rect -1518 -18882 -1508 -18804
rect -1456 -18882 -1446 -18804
rect -1042 -18882 -1032 -18804
rect -980 -18882 -970 -18804
rect -3727 -19016 -802 -18914
rect -3356 -19364 -2226 -19316
rect -2046 -19356 -918 -19316
rect -2046 -19364 -978 -19356
rect -3356 -19536 -3306 -19364
rect -3152 -19472 -3142 -19394
rect -3090 -19472 -3080 -19394
rect -2960 -19472 -2950 -19394
rect -2898 -19472 -2888 -19394
rect -2766 -19472 -2756 -19394
rect -2704 -19472 -2694 -19394
rect -2574 -19472 -2564 -19394
rect -2512 -19472 -2502 -19394
rect -2382 -19472 -2372 -19394
rect -2320 -19472 -2310 -19394
rect -1962 -19472 -1952 -19394
rect -1900 -19472 -1890 -19394
rect -1770 -19472 -1760 -19394
rect -1708 -19472 -1698 -19394
rect -1578 -19472 -1568 -19394
rect -1516 -19472 -1506 -19394
rect -1386 -19472 -1376 -19394
rect -1324 -19472 -1314 -19394
rect -1194 -19472 -1184 -19394
rect -1132 -19472 -1122 -19394
rect -988 -19436 -978 -19364
rect -904 -19436 -894 -19356
rect -3378 -19616 -3368 -19536
rect -3294 -19616 -3284 -19536
rect -3356 -19642 -3306 -19616
rect -3354 -19826 -3306 -19642
rect -2170 -19660 -2102 -19648
rect -3246 -19784 -3236 -19660
rect -3184 -19784 -3174 -19660
rect -3054 -19784 -3044 -19660
rect -2992 -19784 -2982 -19660
rect -2862 -19784 -2852 -19660
rect -2800 -19784 -2790 -19660
rect -2670 -19784 -2660 -19660
rect -2608 -19784 -2598 -19660
rect -2478 -19784 -2468 -19660
rect -2416 -19784 -2406 -19660
rect -2286 -19784 -2276 -19660
rect -2224 -19784 -2214 -19660
rect -2174 -19784 -2164 -19660
rect -2108 -19784 -2098 -19660
rect -2058 -19784 -2048 -19660
rect -1996 -19784 -1986 -19660
rect -1866 -19784 -1856 -19660
rect -1804 -19784 -1794 -19660
rect -1674 -19784 -1664 -19660
rect -1612 -19784 -1602 -19660
rect -1482 -19784 -1472 -19660
rect -1420 -19784 -1410 -19660
rect -1290 -19784 -1280 -19660
rect -1228 -19784 -1218 -19660
rect -1098 -19784 -1088 -19660
rect -1036 -19784 -1026 -19660
rect -2170 -19796 -2102 -19784
rect -966 -19826 -918 -19436
rect -3354 -19874 -2226 -19826
rect -2046 -19874 -918 -19826
<< via1 >>
rect -3088 -15974 -3030 -15854
rect -2772 -15974 -2714 -15854
rect -2456 -15974 -2398 -15854
rect -2162 -15974 -2108 -15854
rect -1872 -15974 -1814 -15854
rect -1556 -15974 -1498 -15854
rect -1240 -15974 -1182 -15854
rect -2930 -16254 -2872 -16134
rect -2614 -16254 -2556 -16134
rect -2298 -16254 -2240 -16134
rect -2030 -16254 -1972 -16134
rect -1714 -16254 -1656 -16134
rect -1398 -16254 -1340 -16134
rect -1962 -16424 -1910 -16372
rect -3560 -17222 -3498 -16990
rect -3082 -17222 -3020 -16990
rect -2606 -17222 -2544 -16990
rect -1750 -17222 -1688 -16990
rect -1274 -17222 -1212 -16990
rect -798 -17222 -736 -16990
rect -3316 -18882 -3264 -18804
rect -2840 -18882 -2788 -18804
rect -2364 -18882 -2312 -18804
rect -1984 -18882 -1932 -18804
rect -1508 -18882 -1456 -18804
rect -1032 -18882 -980 -18804
rect -3142 -19472 -3090 -19394
rect -2950 -19472 -2898 -19394
rect -2756 -19472 -2704 -19394
rect -2564 -19472 -2512 -19394
rect -2372 -19472 -2320 -19394
rect -1952 -19472 -1900 -19394
rect -1760 -19472 -1708 -19394
rect -1568 -19472 -1516 -19394
rect -1376 -19472 -1324 -19394
rect -1184 -19472 -1132 -19394
rect -978 -19436 -904 -19356
rect -3368 -19616 -3294 -19536
rect -3236 -19784 -3184 -19660
rect -3044 -19784 -2992 -19660
rect -2852 -19784 -2800 -19660
rect -2660 -19784 -2608 -19660
rect -2468 -19784 -2416 -19660
rect -2276 -19784 -2224 -19660
rect -2164 -19784 -2108 -19660
rect -2048 -19784 -1996 -19660
rect -1856 -19784 -1804 -19660
rect -1664 -19784 -1612 -19660
rect -1472 -19784 -1420 -19660
rect -1280 -19784 -1228 -19660
rect -1088 -19784 -1036 -19660
<< metal2 >>
rect -3088 -15854 -3030 -15844
rect -2772 -15854 -2714 -15844
rect -2456 -15854 -2398 -15844
rect -2162 -15854 -2108 -15844
rect -1872 -15854 -1814 -15844
rect -1556 -15854 -1498 -15844
rect -1240 -15854 -1182 -15844
rect -3030 -15974 -2772 -15854
rect -2714 -15974 -2456 -15854
rect -2398 -15974 -2162 -15854
rect -2108 -15974 -1872 -15854
rect -1814 -15974 -1556 -15854
rect -1498 -15974 -1240 -15854
rect -1182 -15974 -1118 -15854
rect -3088 -15984 -3030 -15974
rect -2772 -15984 -2714 -15974
rect -2456 -15984 -2398 -15974
rect -2162 -15984 -2108 -15974
rect -1872 -15984 -1814 -15974
rect -1556 -15984 -1498 -15974
rect -1240 -15984 -1182 -15974
rect -2930 -16134 -2872 -16124
rect -2614 -16134 -2556 -16124
rect -2298 -16134 -2240 -16124
rect -3082 -16254 -2930 -16134
rect -2872 -16254 -2614 -16134
rect -2556 -16254 -2298 -16134
rect -2930 -16264 -2872 -16254
rect -2778 -16264 -2556 -16254
rect -2298 -16264 -2240 -16254
rect -2030 -16134 -1972 -16124
rect -1714 -16134 -1656 -16124
rect -1398 -16134 -1340 -16124
rect -1972 -16254 -1714 -16134
rect -1656 -16254 -1398 -16134
rect -1340 -16254 -1188 -16134
rect -2030 -16264 -1972 -16254
rect -1714 -16264 -1520 -16254
rect -1398 -16264 -1340 -16254
rect -3560 -16990 -3498 -16980
rect -3082 -16990 -3020 -16980
rect -2778 -16990 -2680 -16264
rect -2292 -16294 -2244 -16264
rect -2292 -16342 -2090 -16294
rect -2146 -16374 -2090 -16342
rect -1962 -16372 -1910 -16366
rect -2146 -16422 -1962 -16374
rect -1962 -16430 -1910 -16424
rect -2606 -16990 -2544 -16980
rect -3498 -17222 -3082 -16990
rect -3020 -17222 -2606 -16990
rect -3560 -17232 -3498 -17222
rect -3082 -17232 -3020 -17222
rect -2606 -17232 -2544 -17222
rect -1750 -16990 -1688 -16980
rect -1618 -16990 -1520 -16264
rect -1274 -16990 -1212 -16980
rect -798 -16990 -736 -16980
rect -1688 -17222 -1274 -16990
rect -1212 -17222 -798 -16990
rect -1750 -17232 -1688 -17222
rect -1274 -17232 -1212 -17222
rect -798 -17232 -736 -17222
rect -3316 -18804 -3264 -18794
rect -3316 -19054 -3264 -18882
rect -2840 -18804 -2788 -18794
rect -2840 -19054 -2788 -18882
rect -2364 -18804 -2312 -18794
rect -2364 -19054 -2312 -18882
rect -3316 -19140 -2312 -19054
rect -1984 -18804 -1932 -18794
rect -1984 -19054 -1932 -18882
rect -1508 -18804 -1456 -18794
rect -1508 -19054 -1456 -18882
rect -1032 -18804 -980 -18794
rect -1032 -19054 -980 -18882
rect -1984 -19140 -980 -19054
rect -3248 -19248 -2244 -19140
rect -2028 -19248 -1024 -19140
rect -3142 -19394 -3090 -19248
rect -3142 -19482 -3090 -19472
rect -2950 -19394 -2898 -19248
rect -2950 -19482 -2898 -19472
rect -2756 -19394 -2704 -19248
rect -2756 -19482 -2704 -19472
rect -2564 -19394 -2512 -19248
rect -2564 -19482 -2512 -19472
rect -2372 -19394 -2320 -19248
rect -2372 -19482 -2320 -19472
rect -1952 -19394 -1900 -19248
rect -1952 -19482 -1900 -19472
rect -1760 -19394 -1708 -19248
rect -1760 -19482 -1708 -19472
rect -1568 -19394 -1516 -19248
rect -1568 -19482 -1516 -19472
rect -1376 -19394 -1324 -19248
rect -1376 -19482 -1324 -19472
rect -1184 -19394 -1132 -19248
rect -978 -19356 -904 -19346
rect -978 -19446 -904 -19436
rect -1184 -19482 -1132 -19472
rect -3368 -19536 -3294 -19526
rect -3368 -19626 -3294 -19616
rect -3236 -19660 -3184 -19650
rect -3044 -19660 -2992 -19650
rect -2852 -19660 -2800 -19650
rect -2660 -19660 -2608 -19650
rect -2468 -19660 -2416 -19650
rect -2276 -19660 -2224 -19648
rect -2164 -19660 -2108 -19650
rect -2048 -19660 -1996 -19650
rect -1856 -19660 -1804 -19650
rect -1664 -19660 -1612 -19650
rect -1472 -19660 -1420 -19650
rect -1280 -19660 -1228 -19650
rect -1088 -19660 -1036 -19650
rect -3184 -19784 -3044 -19660
rect -2992 -19784 -2852 -19660
rect -2800 -19784 -2660 -19660
rect -2608 -19784 -2468 -19660
rect -2416 -19784 -2276 -19660
rect -2224 -19784 -2164 -19660
rect -2108 -19784 -2048 -19660
rect -1996 -19784 -1856 -19660
rect -1804 -19784 -1664 -19660
rect -1612 -19784 -1472 -19660
rect -1420 -19784 -1280 -19660
rect -1228 -19784 -1088 -19660
rect -3236 -19794 -3184 -19784
rect -3044 -19794 -2992 -19784
rect -2852 -19794 -2800 -19784
rect -2660 -19794 -2608 -19784
rect -2468 -19794 -2416 -19784
rect -2276 -19792 -2224 -19784
rect -2164 -19794 -2108 -19784
rect -2048 -19794 -1996 -19784
rect -1856 -19794 -1804 -19784
rect -1664 -19794 -1612 -19784
rect -1472 -19794 -1420 -19784
rect -1280 -19794 -1228 -19784
rect -1088 -19794 -1036 -19784
<< via2 >>
rect -978 -19436 -904 -19356
rect -3368 -19616 -3294 -19536
<< metal3 >>
rect -988 -19356 -894 -19351
rect -3658 -19436 -978 -19356
rect -904 -19436 -894 -19356
rect -988 -19441 -894 -19436
rect -3378 -19536 -3284 -19531
rect -3658 -19616 -3368 -19536
rect -3294 -19616 -918 -19536
rect -3378 -19621 -3284 -19616
use sky130_fd_pr__nfet_01v8_U85QGS  XM1
timestamp 1644523392
transform 1 0 -2728 0 1 -19595
box -646 -410 646 410
use sky130_fd_pr__pfet_g5v0d10v5_B24TY6  XM5
timestamp 1644523392
transform 1 0 -1606 0 1 -16055
box -624 -496 624 496
use sky130_fd_pr__pfet_g5v0d10v5_B24TY6  XM6
timestamp 1644523392
transform -1 0 -2664 0 1 -16055
box -624 -496 624 496
use sky130_fd_pr__nfet_01v8_U85QGS  sky130_fd_pr__nfet_01v8_U85QGS_0
timestamp 1644523392
transform 1 0 -1542 0 1 -19595
box -646 -410 646 410
use sky130_fd_pr__nfet_05v0_nvt_ARHMTT  sky130_fd_pr__nfet_05v0_nvt_ARHMTT_0
timestamp 1644523392
transform 1 0 -2934 0 1 -17882
box -794 -1258 794 1258
use sky130_fd_pr__nfet_05v0_nvt_ARHMTT  sky130_fd_pr__nfet_05v0_nvt_ARHMTT_1
timestamp 1644523392
transform 1 0 -1364 0 1 -17882
box -794 -1258 794 1258
<< labels >>
rlabel metal3 -3658 -19436 -978 -19356 1 in_n
port 2 n
rlabel metal3 -3658 -19616 -3368 -19536 1 in_p
port 1 n
rlabel metal2 -2778 -17222 -2680 -16134 1 out_n
port 4 n
rlabel metal2 -1618 -17222 -1520 -16134 1 out_p
port 3 n
rlabel metal2 -2108 -19784 -2048 -19660 1 vss_lo
port 6 n
rlabel metal1 -3727 -19016 -3625 -16749 1 vdd_lo
port 7 n
rlabel metal2 -1182 -15974 -1118 -15854 1 vdd_hi
port 5 n
<< end >>
