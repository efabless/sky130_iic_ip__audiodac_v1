magic
tech sky130A
magscale 1 2
timestamp 1645179649
<< metal4 >>
rect 37371 29499 54514 75214
rect 68914 73828 69257 74521
rect 148956 74250 149485 74521
rect 68914 73482 69943 73828
rect 148800 73482 149485 74250
rect 68914 72790 70971 73482
rect 148457 73136 149485 73482
rect 147771 72790 149485 73136
rect 68914 72443 70628 72790
rect 147085 72443 149485 72790
rect 68914 72097 71314 72443
rect 146743 72097 149485 72443
rect 68914 71751 71657 72097
rect 146400 71751 149485 72097
rect 68914 71404 72343 71751
rect 146057 71404 149485 71751
rect 68914 70712 73371 71404
rect 145714 71058 149485 71404
rect 145371 70712 149485 71058
rect 68914 70365 73714 70712
rect 144685 70365 149485 70712
rect 68914 70019 74057 70365
rect 144000 70019 149485 70365
rect 68914 69673 74400 70019
rect 144343 69673 149485 70019
rect 68914 69326 74743 69673
rect 68914 68980 75428 69326
rect 143657 68980 149485 69673
rect 68914 68287 75771 68980
rect 142971 68634 149485 68980
rect 142628 68287 149485 68634
rect 68914 67595 76457 68287
rect 141943 67941 149485 68287
rect 141600 67595 149485 67941
rect 68914 67248 77143 67595
rect 141257 67248 149485 67595
rect 68914 66902 77485 67248
rect 140914 66902 149485 67248
rect 68914 66556 78171 66902
rect 140571 66556 149485 66902
rect 68914 66209 78514 66556
rect 139885 66209 149485 66556
rect 68914 65863 78857 66209
rect 139200 65863 149485 66209
rect 68914 65517 79200 65863
rect 139543 65517 149485 65863
rect 68914 65170 79543 65517
rect 68914 64824 80228 65170
rect 138857 64824 149485 65517
rect 68914 64132 80571 64824
rect 138514 64478 149485 64824
rect 137828 64132 149485 64478
rect 68914 63785 80914 64132
rect 137143 63785 149485 64132
rect 68914 63439 81257 63785
rect 136800 63439 149485 63785
rect 68914 63093 81600 63439
rect 136457 63093 149485 63439
rect 68914 62746 82285 63093
rect 82628 62746 82971 63093
rect 68914 62400 82971 62746
rect 135428 62400 135771 62746
rect 136114 62400 149485 63093
rect 68914 62054 83314 62400
rect 135428 62054 149485 62400
rect 68914 61707 83657 62054
rect 134743 61707 149485 62054
rect 68914 61015 84000 61707
rect 84343 61015 84685 61361
rect 134400 61015 149485 61707
rect 68914 60322 85028 61015
rect 133714 60322 149485 61015
rect 68914 59629 85714 60322
rect 133028 59976 149485 60322
rect 68914 58937 86400 59629
rect 132000 59283 149485 59976
rect 86743 58937 87085 59283
rect 131657 58937 149485 59283
rect 68914 58244 87771 58937
rect 131314 58590 149485 58937
rect 130971 58244 149485 58590
rect 68914 57898 88114 58244
rect 130628 57898 149485 58244
rect 68914 57551 88457 57898
rect 129600 57551 129943 57898
rect 130285 57551 149485 57898
rect 68914 57205 88800 57551
rect 68914 56859 89485 57205
rect 129600 56859 149485 57551
rect 68914 56166 89828 56859
rect 128228 56166 128571 56512
rect 128914 56166 149485 56859
rect 68914 55473 90514 56166
rect 128228 55820 149485 56166
rect 68914 55127 90857 55473
rect 127200 55127 149485 55820
rect 68914 54781 91200 55127
rect 91543 54781 91885 55127
rect 126857 54781 149485 55127
rect 68914 54088 92571 54781
rect 126514 54435 149485 54781
rect 126171 54088 149485 54435
rect 69257 53742 92914 54088
rect 125828 53742 149485 54088
rect 69600 53396 93257 53742
rect 124800 53396 148800 53742
rect 69943 53049 93600 53396
rect 124800 53056 148186 53396
rect 124800 53049 147771 53056
rect 70285 52703 93943 53049
rect 124457 52703 147771 53049
rect 70628 52357 94628 52703
rect 124457 52357 147428 52703
rect 71314 52010 95314 52357
rect 124114 52158 147085 52357
rect 124114 52010 147082 52158
rect 71657 51664 94971 52010
rect 123085 51664 123428 52010
rect 123771 51664 147082 52010
rect 72343 50971 95657 51664
rect 123085 51318 146743 51664
rect 122400 50971 146057 51318
rect 72343 50625 72685 50971
rect 73028 50682 96685 50971
rect 73028 50625 96686 50682
rect 122057 50625 145714 50971
rect 73028 50279 97028 50625
rect 121714 50279 145371 50625
rect 73371 49932 97371 50279
rect 121371 49932 145028 50279
rect 74057 49586 97714 49932
rect 121028 49586 144685 49932
rect 74400 49240 98057 49586
rect 120000 49240 144000 49586
rect 74743 48893 98400 49240
rect 120343 48893 143657 49240
rect 75085 48547 98743 48893
rect 75085 48201 75428 48547
rect 75771 48201 99428 48547
rect 119657 48201 142971 48893
rect 76114 47854 99771 48201
rect 118628 48014 142285 48201
rect 118628 47854 142238 48014
rect 76457 47508 99771 47854
rect 118971 47508 142238 47854
rect 77143 46815 100457 47508
rect 117943 47162 141943 47508
rect 117600 46815 141257 47162
rect 77485 46470 101485 46815
rect 77485 46469 101486 46470
rect 117257 46469 140914 46815
rect 77828 46123 101828 46469
rect 116914 46123 140571 46469
rect 78171 45777 102171 46123
rect 116571 45777 140228 46123
rect 78857 45430 102514 45777
rect 115885 45430 139543 45777
rect 79200 45084 102857 45430
rect 115543 45084 139200 45430
rect 79543 44738 103200 45084
rect 115200 44738 138857 45084
rect 79885 44391 103543 44738
rect 114857 44510 138310 44738
rect 79885 44382 80228 44391
rect 80571 44045 104228 44391
rect 114857 44045 137828 44510
rect 80914 43699 104571 44045
rect 114514 43699 137412 44045
rect 81257 43352 104571 43699
rect 113828 43632 137412 43699
rect 81943 43006 105257 43352
rect 113143 43006 113485 43352
rect 113828 43006 137143 43632
rect 82285 42660 105257 43006
rect 112800 42660 136457 43006
rect 82285 42313 105943 42660
rect 112457 42313 136114 42660
rect 82552 42220 106628 42313
rect 82628 41967 106628 42220
rect 112114 41967 135771 42313
rect 82971 41621 83314 41967
rect 83657 41621 106971 41967
rect 111771 41621 135428 41967
rect 83657 41274 107314 41621
rect 111428 41274 134743 41621
rect 84343 40928 107657 41274
rect 110400 40928 134400 41274
rect 84343 40582 108000 40928
rect 110400 40582 134057 40928
rect 84685 40235 108685 40582
rect 110400 40235 133371 40582
rect 85371 39889 109028 40235
rect 109714 39889 133028 40235
rect 85714 39543 133028 39889
rect 86057 39196 132343 39543
rect 132685 39530 133028 39543
rect 86400 38850 132343 39196
rect 87085 38504 132000 38850
rect 87428 38157 131314 38504
rect 87771 37811 130971 38157
rect 88114 37448 130628 37811
rect 88114 37119 130340 37448
rect 88800 36772 129600 37119
rect 89143 36426 129257 36772
rect 163885 36426 180685 75214
rect 89485 36080 128914 36426
rect 89828 35733 128228 36080
rect 90514 35387 128228 35733
rect 163885 35387 181028 36426
rect 90857 35041 128228 35387
rect 164228 35041 181028 35387
rect 217371 35733 234171 75214
rect 217371 35041 234514 35733
rect 91200 34694 127543 35041
rect 91885 34354 127200 34694
rect 91885 34002 126514 34354
rect 126857 34348 127200 34354
rect 163885 34348 181371 35041
rect 92914 33655 126171 34002
rect 163885 33655 181028 34348
rect 217371 34002 234171 35041
rect 92571 33309 125828 33655
rect 93600 32963 125485 33309
rect 93600 32616 124800 32963
rect 94285 32270 124457 32616
rect 164228 32270 181028 33655
rect 217028 33309 234171 34002
rect 217028 32963 233828 33309
rect 216685 32616 233828 32963
rect 94285 31924 124114 32270
rect 94285 31577 123085 31924
rect 95314 31231 123085 31577
rect 95657 30885 123104 31231
rect 96000 30736 122784 30885
rect 96000 30538 122743 30736
rect 97028 29846 121714 30538
rect 164228 29846 181371 32270
rect 217028 30538 233828 32616
rect 216343 30192 233828 30538
rect 216685 29846 234171 30192
rect 97028 29499 121028 29846
rect 164228 29499 181714 29846
rect 37028 26383 54514 29499
rect 97371 29153 121028 29499
rect 98057 28807 120685 29153
rect 98400 28461 120000 28807
rect 98743 28114 119657 28461
rect 164571 28114 181714 29499
rect 216685 29499 233828 29846
rect 216685 29153 233485 29499
rect 99085 27768 119314 28114
rect 99085 27422 118971 27768
rect 100114 27075 118656 27422
rect 100457 26894 118656 27075
rect 164571 27075 182057 28114
rect 216343 27768 233485 29153
rect 216000 27422 233828 27768
rect 216000 27075 233485 27422
rect 100457 26729 118628 26894
rect 164571 26729 182400 27075
rect 216000 26729 233143 27075
rect 37028 26036 54520 26383
rect 101143 26036 117257 26729
rect 117600 26383 117943 26729
rect 164914 26383 182400 26729
rect 215657 26383 233143 26729
rect 36685 25344 54514 26036
rect 101828 25344 116571 26036
rect 164914 25344 182743 26383
rect 216000 26036 233143 26383
rect 215657 25690 233143 26036
rect 36685 24305 54171 25344
rect 102171 24997 116228 25344
rect 165257 24997 183085 25344
rect 215314 24997 233143 25690
rect 102857 24651 115885 24997
rect 103200 24305 115543 24651
rect 165257 24305 183428 24997
rect 214971 24305 232800 24997
rect 10628 23612 10971 23958
rect 10285 23266 11657 23612
rect 36343 23266 54171 24305
rect 103543 23958 114857 24305
rect 104228 23612 114514 23958
rect 165257 23612 183771 24305
rect 214628 23958 232800 24305
rect 214628 23612 232457 23958
rect 104571 23266 114171 23612
rect 9943 22922 12000 23266
rect 9438 22919 12000 22922
rect 36332 22919 54171 23266
rect 104914 22919 113143 23266
rect 9438 22573 12343 22919
rect 36343 22573 54171 22919
rect 105257 22573 113143 22919
rect 165600 22919 184114 23612
rect 214285 23266 232457 23612
rect 165600 22573 184457 22919
rect 213943 22573 232457 23266
rect 9182 22238 12685 22573
rect 8820 21880 12685 22238
rect 36000 22227 54171 22573
rect 106285 22227 113143 22573
rect 165943 22227 184800 22573
rect 8571 21534 13028 21880
rect 35657 21552 53828 22227
rect 106285 22068 112854 22227
rect 106285 21880 112800 22068
rect 35657 21534 53796 21552
rect 106971 21534 111771 21880
rect 8228 21222 13371 21534
rect 8226 21188 13371 21222
rect 8226 20841 13714 21188
rect 35314 20841 53796 21534
rect 106910 21188 111771 21534
rect 165943 21534 185143 22227
rect 213600 21880 232114 22573
rect 212914 21534 232457 21880
rect 165943 21188 185485 21534
rect 212571 21188 231771 21534
rect 107657 20841 111085 21188
rect 166285 20841 185828 21188
rect 212914 20841 231771 21188
rect 7885 20495 14057 20841
rect 34971 20668 53796 20841
rect 34971 20495 53828 20668
rect 107612 20495 111094 20841
rect 7543 20149 14400 20495
rect 34628 20286 53485 20495
rect 7200 19826 15180 20149
rect 7200 19803 15428 19826
rect 6857 19456 15428 19803
rect 34608 19656 53485 20286
rect 108343 20149 110743 20495
rect 166285 20149 186514 20841
rect 212228 20495 231771 20841
rect 212228 20149 231428 20495
rect 108343 19803 110057 20149
rect 166628 19803 186857 20149
rect 211200 19803 231428 20149
rect 34628 19456 53485 19656
rect 108685 19456 109714 19803
rect 166628 19456 187200 19803
rect 211543 19456 231428 19803
rect 6514 19110 16114 19456
rect 33943 19110 53485 19456
rect 166628 19116 187885 19456
rect 166628 19110 187890 19116
rect 210514 19110 231085 19456
rect 6044 18924 16457 19110
rect 5828 18764 16457 18924
rect 33600 18764 53143 19110
rect 5828 18417 16800 18764
rect 5485 18071 17143 18417
rect 33272 18296 53143 18764
rect 166971 18417 188571 19110
rect 210857 18764 231085 19110
rect 209828 18417 230743 18764
rect 33257 18071 53143 18296
rect 108343 18071 109028 18072
rect 167314 18071 189257 18417
rect 209143 18071 230743 18417
rect 5485 17725 17828 18071
rect 32228 17784 52800 18071
rect 5143 17378 18857 17725
rect 32126 17378 52800 17784
rect 4800 17032 19200 17378
rect 31543 17032 52800 17378
rect 4457 16686 19885 17032
rect 30514 16686 30857 16694
rect 31200 16686 52457 17032
rect 4114 16339 21257 16686
rect 28800 16339 29143 16340
rect 29828 16339 52457 16686
rect 3771 15993 21943 16339
rect 22285 15993 22971 16339
rect 28457 15993 52482 16339
rect 3771 15864 52114 15993
rect 3280 15300 52114 15864
rect 2743 14954 52114 15300
rect 3085 14608 51771 14954
rect 2400 14261 51771 14608
rect 1714 14236 2057 14261
rect 2400 14236 51428 14261
rect 1714 13915 51428 14236
rect 1714 13569 51085 13915
rect 1371 13222 51085 13569
rect 1028 12876 51090 13222
rect 685 12530 50743 12876
rect 343 12183 50743 12530
rect 338 11837 50400 12183
rect 685 11491 50057 11837
rect 1028 11144 50057 11491
rect 1028 10798 49714 11144
rect 1371 10472 49714 10798
rect 1371 10452 49226 10472
rect 1714 10106 49028 10452
rect 2057 9759 49028 10106
rect 2400 9413 48685 9759
rect 2743 9067 48343 9413
rect 3085 8720 48343 9067
rect 3428 8374 48000 8720
rect 3771 8028 47657 8374
rect 3966 8020 47314 8028
rect 4457 7681 47314 8020
rect 4457 7335 46971 7681
rect 5143 6989 46628 7335
rect 5485 6642 46285 6989
rect 5828 6296 45943 6642
rect 6171 5950 45600 6296
rect 6320 5922 45257 5950
rect 7200 5646 45257 5922
rect 7200 5257 44571 5646
rect 44914 5603 45257 5646
rect 7885 4911 44571 5257
rect 8571 4564 43543 4911
rect 9257 4218 42857 4564
rect 9600 3872 42514 4218
rect 10628 3525 41828 3872
rect 10971 3179 41143 3525
rect 11657 2833 40457 3179
rect 12685 2486 39771 2833
rect 40114 2784 40457 2833
rect 13371 2140 38400 2486
rect 38743 2450 39085 2486
rect 14400 1794 37714 2140
rect 15428 1448 37028 1794
rect 16800 1101 35657 1448
rect 68914 1101 149485 18071
rect 167314 17725 189600 18071
rect 208800 17725 230743 18071
rect 167657 17378 189600 17725
rect 207771 17378 230400 17725
rect 167657 17032 190971 17378
rect 207428 17032 230400 17378
rect 168000 16686 192000 17032
rect 206400 16686 230057 17032
rect 168000 16339 192685 16686
rect 205371 16339 230057 16686
rect 168343 15993 194400 16339
rect 204000 15993 229714 16339
rect 168343 15647 196114 15993
rect 202285 15647 229714 15993
rect 168685 14954 229371 15647
rect 169028 14261 229028 14954
rect 169371 14026 229028 14261
rect 169371 13915 228343 14026
rect 228685 13915 229028 14026
rect 170057 13569 228343 13915
rect 170057 13222 228324 13569
rect 170057 12876 228343 13222
rect 170400 12183 227657 12876
rect 170743 11837 227314 12183
rect 171085 11491 226971 11837
rect 171085 11144 226628 11491
rect 171085 10798 171428 11144
rect 171771 10798 226285 11144
rect 172114 10452 225943 10798
rect 172800 10106 225943 10452
rect 172800 9413 225600 10106
rect 173143 9067 225257 9413
rect 173485 8720 224914 9067
rect 173828 8374 224228 8720
rect 174514 8028 223885 8374
rect 174857 7681 223200 8028
rect 174857 7335 175200 7681
rect 175543 7335 222857 7681
rect 174857 6989 222514 7335
rect 176228 6642 222171 6989
rect 176228 6296 221828 6642
rect 176571 5950 221143 6296
rect 177257 5603 220800 5950
rect 177600 5257 220114 5603
rect 178285 4911 220114 5257
rect 178971 4564 219085 4911
rect 179657 4218 218057 4564
rect 180000 3872 217714 4218
rect 181028 3525 217028 3872
rect 181714 3179 216343 3525
rect 182057 2833 215657 3179
rect 183085 2486 214628 2833
rect 184114 2140 213600 2486
rect 185143 1794 212571 2140
rect 213257 1794 213600 2140
rect 186171 1448 186514 1794
rect 186857 1448 210857 1794
rect 211200 1448 211543 1794
rect 187543 1101 210171 1448
rect 18171 755 34285 1101
rect 188914 755 189257 1101
rect 189600 755 208800 1101
rect 20228 409 32228 755
rect 191314 409 206400 755
rect 20571 372 20914 409
rect 22971 62 29485 409
rect 31543 392 31885 409
rect 193371 62 202971 409
rect 203314 62 204343 409
rect 24343 0 24685 62
rect 27771 0 28114 62
<< end >>
